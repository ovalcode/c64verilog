`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05.07.2017 15:35:00
// Design Name: 
// Module Name: test
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module test(
  input clk,
  output [7:0] led
    );
    
    
    
    
    //wire [7:0] DO;
//    reg clk = 0;
    reg [15:0] addr = 16'h2461;
//    reg reset = 1;
    reg EN = 0;
    
    wire [7:0] DATA_OUT_BLOCK_0;
    wire [7:0] DATA_OUT_BLOCK_1;
    wire [7:0] DATA_OUT_BLOCK_2;
    wire [7:0] DATA_OUT_BLOCK_3;
    wire [7:0] DATA_OUT_BLOCK_4;
    wire clk_out;
    wire nc_wire;
    reg [7:0] combined_data_out;
    reg [24:0] clk_counter = 0;
    
    
clk_wiz_0 clk_gen 
         (
          // Clock out ports
          clk_out,
          // Status and control signals
          0,
          nc_wire,
         // Clock in ports
          clk
         );


    assign led = combined_data_out;
/*    initial begin
      #1000000;
      EN <= 1;
      reset <= 0;
      #100;
      //EN <= 0;
    end*/
    
 
   BRAM_SINGLE_MACRO #(
       .BRAM_SIZE("36Kb"), // Target BRAM, "18Kb" or "36Kb" 
       .DEVICE("7SERIES"), // Target Device: "7SERIES" 
       .DO_REG(0), // Optional output register (0 or 1)
       .INIT(36'h000000000), // Initial values on output port
       .INIT_FILE ("NONE"),
       .WRITE_WIDTH(8), // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
       .READ_WIDTH(8),  // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
       .SRVAL(36'h000000000), // Set/Reset value for port output
       .WRITE_MODE("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE" 
       .INIT_00(256'hA89FA9A4AC05B080ABBEABA4A8F7AD1DA741A83043495341424D4243E37BE394),
       .INIT_01(256'hAA9FAA7FB823B3B2E164E155E167B82CA94AA82EA93AA8D1A882A81CA927A870),
       .INIT_02(256'hBF71B39EB37D0310BC58BCCCBC39A641AB7AE1C6E1BDE129AA85A65DA69BA856),
       .INIT_03(256'hB737B72CB700B6ECB78BB7ADB465B77CB80DE30EE2B4E26BE264BFEDB9EAE097),
       .INIT_04(256'h4E45B01564AED35ABFB37DAFE546AFE850BF7A7FBB117BBA2A7BB85279B86979),
       .INIT_05(256'h454CC4414552CD4944D455504E49A35455504E49C1544144D458454ED24F46C4),
       .INIT_06(256'h53CD4552CE5255544552C255534F47C5524F54534552C649CE5552CF544F47D4),
       .INIT_07(256'h5250C54B4F50C64544D94649524556C5564153C4414F4CD4494157CE4FD04F54),
       .INIT_08(256'h4C43CE45504FD35953C44D43D24C43D453494CD44E4F43D44E495250A3544E49),
       .INIT_09(256'hD0455453D44F4ECE454854A8435053CE46CF54A8424154D7454ED44547C5534F),
       .INIT_0A(256'h53D34F50C55246D25355D34241D44E49CE4753BCBDBED24FC44E41DEAFAAADAB),
       .INIT_0B(256'h5453CE454CCB454550CE5441CE4154CE4953D34F43D05845C74F4CC44E52D251),
       .INIT_0C(256'h4F5400CF47A444494DA45448474952A45446454CA4524843C35341CC4156A452),
       .INIT_0D(256'h504F20544F4E20454C4946CE45504F20454C4946D3454C494620594E414D204F),
       .INIT_0E(256'h455345525020544F4E20454349564544C44E554F4620544F4E20454C4946CE45),
       .INIT_0F(256'h4DC54C49462054555054554F20544F4EC54C4946205455504E4920544F4ED44E),
       .INIT_10(256'h4E20454349564544204C4147454C4C49C54D414E20454C494620474E49535349),
       .INIT_11(256'h5255544552D841544E5953D24F462054554F48544957205458454ED245424D55),
       .INIT_12(256'h4147454C4C49C154414420464F2054554FC255534F472054554F48544957204E),
       .INIT_13(256'h55D9524F4D454D20464F2054554FD74F4C465245564FD95449544E415551204C),
       .INIT_14(256'h444552D4504952435342555320444142D44E454D45544154532044274645444E),
       .INIT_15(256'h4147454C4C49CF52455A205942204E4F495349564944D9415252412044274D49),
       .INIT_16(256'h204F4F5420474E49525453C84354414D53494D2045505954D44345524944204C),
       .INIT_17(256'hD8454C504D4F43204F4F5420414C554D524F46C154414420454C4946C74E4F4C),
       .INIT_18(256'h4556CE4F4954434E55462044274645444E55C5554E49544E4F432054274E4143),
       .INIT_19(256'hA23BA235A225A210A1FFA1F0A1E2A1D0A1C2A1B5A1ACA19EC4414F4CD9464952),
       .INIT_1A(256'hA31EA30EA300A2EDA2E4A2D5A2C8A2BAA2AAA29DA290A27FA272A26AA25AA24F),
       .INIT_1B(256'h0A0D2E59444145520A0D00204E492000524F5252452020000D4B4F0DA383A324),
       .INIT_1C(256'hBD49850102BD0AD04AA521D081C90101BDE8E8E8E8BAA0004B414552420A0D00),
       .INIT_1D(256'h3832843185A4082060D8D0AA1269188A07F00102DD49A507D00103DD4A850103),
       .INIT_1E(256'h22E558A5385BC603B05A8522E5385AA523F098E8AA60E55BA5A822855FE55AA5),
       .INIT_1F(256'h35B03E690A60F2D0CA59C65BC658915AB1F9D08858915AB1049059C608B05885),
       .INIT_20(256'hA2B52620FA10CA57B5489809A248229033C504D0289034C4602E9022E4BA2285),
       .INIT_21(256'hA326BDAA0A8A03006C10A26001B033C505D0069034C468A868FA30E8619568F7),
       .INIT_22(256'h68C8AB47207F294822B100A0AB4520AAD720138500A9FFCC202385A327BD2285),
       .INIT_23(256'hFF902080A9AB1E20A3A076A9BDC22003F0C83AA4AB1E20A3A069A9A67A20F410),
       .INIT_24(256'h20A96B20A7E14CA5792006903A86FFA2F0F0AA0073207B847A86A5602003026C),
       .INIT_25(256'h852D65185FF1885FA5258560A522852DA523855FB101A04490A613200B84A579),
       .INIT_26(256'hB11823C6039022651825C6E803B0A82DE55FA538AA60E52E85FF692EA524852D),
       .INIT_27(256'h850B655A852DA51888F00200ADA53320A65920F2D0CA25E623E6F9D0C8249122),
       .INIT_28(256'hA42E842D8532A431A501FF8C01FE8D15A414A5A3B8205984C801905B842EA458),
       .INIT_29(256'h22B101A018238422852CA42BA5A4804CA53320A65920F810885F9101FCB9880B),
       .INIT_2A(256'h60DD90238522862291C8006923A5229100A0AA226598C8FBD022B1C804A01DF0),
       .INIT_2B(256'h04A07AA603046CAACA4CA4374C17A2F19059E0E802009D0DF00DC9E1122000A2),
       .INIT_2C(256'h04D03FC92D700F2456F022C9088537F020C9F4D0E83EF0FFC907100200BD0F84),
       .INIT_2D(256'hF0A09EF9380200BDE8C8CA7A86880B8400A071841D903CC9049030C925D099A9),
       .INIT_2E(256'hE9380F8502D049C904F03AE93836F001FBB901FB99C8E871A40B0530D080C9F5),
       .INIT_2F(256'hB9FA10A09DB9C80BE67AA6F0D0E801FB99C8DBF008C5DFF00200BD08859FD055),
       .INIT_30(256'hF05FB160865F8501A02CA62BA5607A85FFA97BC601FD99BE100200BDB4D0A09E),
       .INIT_31(256'hD7B05FB188AA5FB1880AF00C905FD18814A509D08803F018905FD115A5C8C81F),
       .INIT_32(256'h2DD000A9A68E202E8500692CA52D850269182BA52B91C82B91A800A9FDD06018),
       .INIT_33(256'hA868168619A2A81D203284318530842F852EA42DA53484338538A437A5FFE720),
       .INIT_34(256'h04F00690607B85FF692CA57A85FF692BA5186010853E8500A94898489AFAA268),
       .INIT_35(256'h0514A5686886D0A96B200073208ED0ABC90CF0007920A61320A96B20E9D0ABC9),
       .INIT_36(256'h15C55FB1C8AA5FB1C8AAD720A82C2043F05FB10F8401A015851485FFA906D015),
       .INIT_37(256'h0F85FF490FA506D022C9AB47207F2949A420A9BDCD2049842CB002F014E404D0),
       .INIT_38(256'hD3F0FFC9D71003066CE3864CB5D060855F865FB1C8AA5FB1A810D05FB111F0C8),
       .INIT_39(256'hAB4720B230A09EB9C8F530FA10A09EB9C808F0CAFFA04984AA7FE938CF300F24),
       .INIT_3A(256'h659818A90620A3FB2009A968689AAA0F698A05D0A38A20A9A520108580A9F5D0),
       .INIT_3B(256'h628562257F0966A5AD8A20AD8D20AEFF20A4A94839A5483AA54800697BA5487A),
       .INIT_3C(256'h20AD8A2000732006D0A9C9007920BBA220B9A0BCA9AE434C23842285A7A08BA9),
       .INIT_3D(256'h00A03E843D8504F0EA02C07BA47AA5A82C204881A94849A5484AA5AE3820BC2B),
       .INIT_3E(256'hE602907A857A65983A857AB1C839857AB1C8A84B4C03D0187AB102A043D07AB1),
       .INIT_3F(256'hA00CB948A00DB9A80A17B023C9119080E93CF0A7AE4CA7ED2000732003086C7B),
       .INIT_40(256'h2BA538A8A04CAEFF20A4A9007320F9D04BC9AF084CD6F03AC9A9A54C00734C48),
       .INIT_41(256'h843D850CF0E83AA67BA47AA53CD01801B0FFE12060428441858801B02CA401E9),
       .INIT_42(256'h4C03D03EA41AA217D0E3864CA4694C0390A3A081A968683C843B853AA439A53E),
       .INIT_43(256'hA66020A6594C03D028FF902000A908603A8439853CA43BA57B847A853DA5A437),
       .INIT_44(256'hA7AE4CA8A020007920488DA94839A5483AA5487AA5487BA5A3FB2003A9A8974C),
       .INIT_45(256'h2CA62BA504B0E807907BA67A6538980BB015E53AA514E539A538A90920A96B20),
       .INIT_46(256'h0BF08DC99AA38A204A85FFA9FDD0607B8500E960A57A8501E95FA51E90A61720),
       .INIT_47(256'h857A651898A906207B85687A85683A856839856868AF084CA4374C11A22C0CA2),
       .INIT_48(256'hF008C5E8F07AB10886078507A608A5088400A0078600A22C3AA2607BE602907A),
       .INIT_49(256'hBBF0A9092005D061A5AEFF20A7A905F089C9007920AD9E20E9F0F3D022C9C8E4),
       .INIT_4A(256'h20A7EF4C6804D065C691D089C904F08DC948B79E20A7ED4CA8A04C03B0007920),
       .INIT_4B(256'hA5D4B019C9228515A507852FE9F7B01586148600A26068EEF02CC9A96B200073),
       .INIT_4C(256'h2015E602901485076514A5152614061585156522A51485146522260A22260A14),
       .INIT_4D(256'hD0AD90202A68AD9E20480DA5480EA5AEFF20B2A94A844985B08B20A9714C0073),
       .INIT_4E(256'h4CD0BFC04AA468BBD04C60499165A5C8499164A500A0B1BF20BC1B2012106818),
       .INIT_4F(256'hAABC0C20AA1D2071A471E6BAE220AA1D2071846684618400A03DD006C9B6A620),
       .INIT_50(256'h2022B1FFDB4C65A563A464A6BC9B20BAE220DFD006C0C871A4BAED208AE805F0),
       .INIT_51(256'hC465A40E9033C564B18807D0179034C564B102A0BD7E4C2FE9B2484C03900080),
       .INIT_52(256'h846F8551A450A5B4752064B100A0AA684C65A464A507B02DC564A50DD008902E),
       .INIT_53(256'h60499150B1C8499150B1C8499150B100A0B6DB205184508500A061A9B67A2070),
       .INIT_54(256'h007920AB2120AAA04C28E11820138608AEFF202CA905F0B79E20ABB54CAA8620),
       .INIT_55(256'h20BDDD20DE300D24AD9E205EF03BC937F02CC94BF018A6C950F0A3C943F035F0),
       .INIT_56(256'h05101324AB47200DA910D013A501A0FFA202009D00A9D3D0AB3B20AB2120B487),
       .INIT_57(256'h200984FFF020380816D00169FF49FCB00AE93898FFF0203860FF49AB47200AA9),
       .INIT_58(256'h8720F2D0AB3B20AAA24C00732006D0CAE8AA059009E58A06902859D029C9B79B),
       .INIT_59(256'hA903F013A5AB284CAAE520F3D00DC9C8AB472022B1BCF0CAE800A0AAB6A620B4),
       .INIT_5A(256'h4C3A84398540A43FA504D0FFA0043011F011A560FF29E10C203FA92C1DA92C20),
       .INIT_5B(256'h23C9B3A620607B847A853EA43DA5AB1E20ADA00CA9A4374C18A205F013A5AF08),
       .INIT_5C(256'hAC0F2040A902018D00A902A001A2E11E201386AEFF202CA9B79E2000732010D0),
       .INIT_5D(256'hC960138600A2FFCC2013A5ABCE20E11E201386AEFF202CA9B79E206013D013A6),
       .INIT_5E(256'hFFB7200DF013A5ABF92001FF8D2CA9B3A620AB2120AEFF203BA9AEBD200BD022),
       .INIT_5F(256'hAB452006D013A5A8FB4CA90620E3D013A51ED00200ADA8F84CABB52006F00229),
       .INIT_60(256'h7BA47AA54A844985B08B2044844386118500A92C98A942A441A6A5604CAB3B20),
       .INIT_61(256'hD001A0FFA202008DE124200C50112420D00079207B847A8644A443A64C844B85),
       .INIT_62(256'hA97A86E80950112431100D240073207B847A86ABF920AB452003D013A575300C),
       .INIT_63(256'hB48D20C8019000697BA47AA50885182CA907853AA907F022C907850CF0078500),
       .INIT_64(256'hA47AA5AB4D4C03F02CC907F0007920A9C2200EA5BCF320AC914CA9DA20B7E220),
       .INIT_65(256'hA212D0AAC8A90620AC154CAEFD202DF00079207B847A854CA44BA5448443857B),
       .INIT_66(256'hA5AC514CDCD083E0AA007920A8FB204085C87AB1C83F857AB1C86CF07AB1C80D),
       .INIT_67(256'h5458453F60AB1E4CACA0FCA907D013A50BF043B100A0A8274C031011A644A443),
       .INIT_68(256'h04D0000D5452415453204D4F5246204F4445523F000D4445524F4E4749204152),
       .INIT_69(256'h6824850669480469188A9AA4374C0AA205F0A38A204A844985B08B2003F000A0),
       .INIT_6A(256'hF00109FD38BABC5D2001A0BBD020B867204AA449A566850109BDBABBA22001A0),
       .INIT_6B(256'h0079209AAA11698AA7AE4C7B850111BD7A850112BD3A850110BD3985010FBD17),
       .INIT_6C(256'h7AA6A4374C16A2FDB06003B003300D24382418AD9E20AD2420007320F1D02CC9),
       .INIT_6D(256'h1790B1E9380079204D8500A9AE8320A3FB2001A9488A482400A27AC67BC602D0),
       .INIT_6E(256'h9007697BB02CD04DA6ADBB4C0073204D8561904DC54D4501492A01C913B003C9),
       .INIT_6F(256'h4BA468AE202048AD8D2067B0A080D968A822650A2285FF69B63D4C03D00D6577),
       .INIT_70(256'hD99048B0A080D9D7D04D851BA07AC67BC602D07AA62A8A0D465FD056F0AA1710),
       .INIT_71(256'h856822E6228568A8A080BE66A5AF084CADA94C4DA5AE332048A081B948A082B9),
       .INIT_72(256'hF064C923F068FFA000226C4861A54862A54863A54864A54865A5BC1B20489823),
       .INIT_73(256'h6F8566456E85686D85686C85686B85686A856869856812854A684B84AD8D2003),
       .INIT_74(256'hA8A90FD0FFC9AF284C0390B11320BCF34C03B00073200D8500A9030A6C6061A5),
       .INIT_75(256'hA47AA50FD022C9D1F0AAC958F0ABC9DEF02EC9A1DA0F498200734CBBA220AEA0),
       .INIT_76(256'hFF4964A5A8FF4965A5B1BF203BD018A013D0A8C9B7E24CB48720C8019000697B),
       .INIT_77(256'hA02CA92C28A92C29A9AD9E20AEFA20AFA74C0390B4C9B3F44C03D0A5C9B3914C),
       .INIT_78(256'hA90890A0E965A500E964A538ADFA4C686815A0A4374C0BA200734C03D07AD100),
       .INIT_79(256'h1C90AF1420708500A926F00DA546A445A665846485B08B206065E5E3A964E5A2),
       .INIT_7A(256'h100E2460B46F4CBE682024A05D8406A07184885E84AF842014D0C9C018D054E0),
       .INIT_7B(256'hA298AF842025D049C01BD054E02D90AF1420B3914C8AA864B1C8AA64B100A00D),
       .INIT_7C(256'hBC3C4CFFB72006D054C00AD053E060628400A0658563846486FFDE20BC4F4CA0),
       .INIT_7D(256'hA5AA68AD8F20AEFD20AD9E20AEFA2020908FE0007320AA480ABBA24C65A464A5),
       .INIT_7E(256'h56859FEBB955859FEAB9A868AEF120AFD64C488AA868B79E20488A4864A54865),
       .INIT_7F(256'h20BBFC2008850B4565A507850B4564A5B1BF200B8400A02CFFA0AD8D4C005420),
       
       // The next set of INITP_xx are for the parity bits
       .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
       
       // The next set of INIT_xx are valid when configured as 36Kb
       .INITP_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0F(256'h0000000000000000000000000000000000000000000000000000000000000000)
    ) BRAM_SINGLE_MACRO_inst_BLOCK_0 (
       .DO(DATA_OUT_BLOCK_0),       // Output data, width defined by READ_WIDTH parameter
       .ADDR(addr[11:0]),   // Input address, width defined by read/write port depth
       .CLK(clk_counter[24]),     // 1-bit input clock
       .DI(0),       // Input data port, width defined by WRITE_WIDTH parameter
       .EN(1),       // 1-bit input RAM enable
       .REGCE(0), // 1-bit input output register enable
       .RST(0),     // 1-bit input reset
       .WE(8'h00)        // Input write enable, width defined by write port depth
    );
 
 
 //===============================================================================================
 
    BRAM_SINGLE_MACRO #(
       .BRAM_SIZE("36Kb"), // Target BRAM, "18Kb" or "36Kb" 
       .DEVICE("7SERIES"), // Target Device: "7SERIES" 
       .DO_REG(0), // Optional output register (0 or 1)
       .INIT(36'h000000000), // Initial values on output port
       .INIT_FILE ("NONE"),
       .WRITE_WIDTH(8), // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
       .READ_WIDTH(8),  // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
       .SRVAL(36'h000000000), // Set/Reset value for port output
       .WRITE_MODE("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE" 
       .INIT_00(256'h257F096EA513B0AD9020B3914C0B4507250B4564A5A80B4508250B4565A5B1BF),
       .INIT_01(256'hA46CA5638462866185B6A6204DC60D8500A9B0614CAABC5B2000A069A96A856A),
       .INIT_02(256'hA607D0CAC8E8FFA06685FFA961A6049001A908F061E538AA6D846C86B6AA206D),
       .INIT_03(256'hFD20BC3C4CFFA902F012252A8AE801A202B0FFA2EFF062D16CB10C90180F3066),
       .INIT_04(256'hA2AF084C03B0B1132000792045850C8600792000A260F4D0007920B09020AAAE),
       .INIT_05(256'hFFA906D024C9F6B0B11320FB90007320AA0B90B1132005900073200E860D8600),
       .INIT_06(256'h1005384686007320AA80098A458545050E8580A9D0D010A513D025C910D00D85),
       .INIT_07(256'hD05FD145A522F02FC504D030E45F8560862EA62DA5108400A0B1D14C03D028E9),
       .INIT_08(256'hC9486860A5E9385BE9059041C9DCD0E8E19007695FA518887DF05FD1C846A508),
       .INIT_09(256'hC004D053C9AF084C03D049C0EFF0C9C00BD054C946A445A560BFA013A905D02A),
       .INIT_0A(256'hA3B82059845885C801900769185B845A8532A431A560845F8530A42FA5F5F054),
       .INIT_0B(256'hC85F91C85F91C85F91C800A95F9146A5C85F9145A500A030842F85C859A458A5),
       .INIT_0C(256'hC8019060A45F6505690A0BA56048844785C8019060A40269185FA55F91C85F91),
       .INIT_0D(256'hA50D3066A5AD8D20AD9E200073206065A464A5B1BF2000000080906059845885),
       .INIT_0E(256'h4846A5489800A0480DA5480E050CA5BC9B4C7AD0BC5B20B1A0A5A9099090C961),
       .INIT_0F(256'h019D65A501029D64A5480101BD480102BDBAA868468568458568B1B2204845A5),
       .INIT_10(256'h60855F8630A52FA60C857F290E85680D8568AEF7200B84D2F02CC9007920C801),
       .INIT_11(256'hB1C8AA5F65185FB1C816F05FD146A506D045C5C85FB100A039F031E404D032C5),
       .INIT_12(256'hEA4CE7D05FD104A00BA5B19420F7D00CA513A2A4374C0EA22C12A2D79060655F),
       .INIT_13(256'hA57186CACA02105F9146A5C8CA01105F9145A505A2728400A0A40820B19420B2),
       .INIT_14(256'hB34C205F918AC85F91C8006968AA0169186808500C2400A90BA25F91C8C8C80B),
       .INIT_15(256'h32843185A4082052F0C8039058658AA859855DB05965DCD00BC622A472857186),
       .INIT_16(256'h32A55F9102A05FE531A53859E6F5D072C659C6FBD058918805F071A472E600A9),
       .INIT_17(256'h0E905FD16585686485AA68C87285718500A90B855FB1C862D00CA55F9160E5C8),
       .INIT_18(256'h22A498AA64658AB34C200AF018710572A5C8A4354CB2454C07905FD18AC806D0),
       .INIT_19(256'h658AB3552000A92886CACA021046A5CA011045A505A27285CAD00BC671866565),
       .INIT_1A(256'h8A00A000A25D8510A929855FB18828855FB122846047A5A84885596598478558),
       .INIT_1B(256'hF00DA560E3D05DC693B0A8296598AA28658A180B9072267106A4B0A82A98AA0A),
       .INIT_1C(256'h2038BC444C90A2638462850D8600A232E534A5A831E533A538B52620B6A62003),
       .INIT_1D(256'h108580A9AEFA20B3A620B3E120A4374C1BA22C15A2A0D0E83AA6EBF000A9FFF0),
       .INIT_1E(256'h4F4CA8F820487AA5487BA54847A54848A548AEFF20B2A9AEF720AD8D20B08B20),
       .INIT_1F(256'hAEF120484EA5484FA5B3E120AD8D4C4F844E85B0922010858009AEFF20A5A9B4),
       .INIT_20(256'h48A4FA10884847B1C8488599F04EB1C8AA47854EB102A04F85684E8568AD8D20),
       .INIT_21(256'h85684E8568AD8A204847A54848A57B854EB1C87A854EB1487AA5487BA5BBD420),
       .INIT_22(256'h4E91C8684E91C8684E91C8684E916800A07B85687A8568AF084C03F00079204F),
       .INIT_23(256'hB4F4205184508665A464A612F000A0FFA96868BDDF2000A0AD8D20604E91C868),
       .INIT_24(256'h04F007C50CF06FB1C8FFA06384628570846F850886078622A260618563846286),
       .INIT_25(256'h980BD002C904F070A57286E8019070A671856F659861841801F022C9F3D008C5),
       .INIT_26(256'h9563A5019562A5009561A5A4374C19A205D022E016A6B6882070A46FA6B47520),
       .INIT_27(256'h01B034A4336538FF49480F46601686E8E8E817860D848870846584648600A002),
       .INIT_28(256'hA9B52620B6300FA510A26068AA36843585348433850B9031C504D0119032C488),
       .INIT_29(256'h00A219A960865F8532A631A54E844F8400A03485338638A537A6D0D0680F8580),
       .INIT_2A(256'hF02FC504D030E4238622852EA62DA5538507A9F7F0B5C72005F016C523862285),
       .INIT_2B(256'h862285B6064C03D031C507D032E459A658A5538503A959865885F3F0B5BD2005),
       .INIT_2C(256'hB1C8D0308AD310285985596522B1C85885586522B1C80822B1C8AA22B100A023),
       .INIT_2D(256'h3022B1F3F0B5C720BAF058C504D059E423A623E602902285226505690A00A022),
       .INIT_2E(256'h169060C51AB033E41ED0069034C522B1C8AA22B1C82BF022B1C8301022B1C835),
       .INIT_2F(256'hE60290228522651853A5558553A54F864E8523A622A560855F8610905FE404D0),
       .INIT_30(256'h5B85006960A55A855F654EB15585A84A042955A5F5F04E054FA56000A023A623),
       .INIT_31(256'h4865A5B52A4C4E91C859A559E6AA4E9158A5C855A4A3BF205986588534A633A5),
       .INIT_32(256'hB47520A4374C17A205906471186FB100A07085686F8568AD8F20AE83204864A5),
       .INIT_33(256'hC8486FB100A0ADB84CB4CA20B6AA2070A46FA5B68C20B6AA2051A450A5B67A20),
       .INIT_34(256'h0290358535651868F8D098359122B188480AF0A82384228668A86FB1C8AA6FB1),
       .INIT_35(256'h68A822B1C8AA22B1C84822B100A008B6DB202384228565A464A5AD8F206036E6),
       .INIT_36(256'hC50CD018C460238422866834E602903385336518480BD033E40FD034C413D028),
       .INIT_37(256'hB4CA4C6868629100A068B47D2001A9488AB7A1206000A0178503E9168508D017),
       .INIT_38(256'h8522651868A868B6AA2051A450A5B47D20488A4898AA50B104909850D1B76120),
       .INIT_39(256'h29C90079206585FFA9B7064CFF4950F118B76120B4CA4CB68C209823E6029022),
       .INIT_3A(256'hB065A5B19065C5FF49B6B050F100A218488ACA4BF0B76120B79E20AEFD2006F0),
       .INIT_3B(256'h4CB78220608A00A048984855A5518568508568AA686868558568A868AEF720AD),
       .INIT_3C(256'h8A20007320B2484CB3A24CA822B100A008F0B7822060A80D8600A2B6A320B3A2),
       .INIT_3D(256'h8622A6728471867BA47AA6B8F74C03D0B7822000794C65A6F0D064A6B1B820AD),
       .INIT_3E(256'h00A068BCF3200079202491984824B100A02586E801907B8623A624852265187A),
       .INIT_3F(256'hB091C961A59D3066A5B79E4CAEFD20B7F720AD8A20607B847A8672A471A62491),
       .INIT_40(256'h8568148568A814B100A0B7F7204814A54815A5601585148465A464A5BC9B2097),
       .INIT_41(256'h00A04A86B7F12003F000792000A24986B7EB2060149100A08AB7EB20B3A24C15),
       .INIT_42(256'h4C61A56F856E456685FF4966A5BA8C20B8674CBFA011A960F8F049254A4514B1),
       .INIT_43(256'h9024F061E538CEF0A869A569A2568670A6BBFC4C03D0BA8C203C90B99920B86A),
       .INIT_44(256'h015670A5A8C730F9C9708400A004D061A2568400A00069FF4966846EA4618412),
       .INIT_45(256'h0003B9658504F50004B970855665FF493869A002F069E061A057106F24B9B020),
       .INIT_46(256'hA64AD062A6189800A0B9472003B0628501F50001B9638502F50002B9648503F5),
       .INIT_47(256'h5665606685618500A9E4D020C908697084658670A6648665A6638664A6628663),
       .INIT_48(256'h060169B9364C62856A6562A563856B6563A564856C6564A565856D6565A57085),
       .INIT_49(256'h6366626642F061E60E9061850169FF49C7B061E538F210622663266426652670),
       .INIT_4A(256'hA56485FF4964A56385FF4963A56285FF4962A56685FF4966A560706665666466),
       .INIT_4B(256'h0FA26062E602D063E606D064E60AD065E60ED070E67085FF4970A56585FF4965),
       .INIT_4C(256'hE9E6F0E8300869019468A4029401B4039402B4049403B4708404B425A2A4374C),
       .INIT_4D(256'h000000816018ECD0C86A0476037602760176017601F60290011614B070A5A808),
       .INIT_4E(256'h34F304358134F3043580203BAA38821693387680640B9B138079CB565E7F0300),
       .INIT_4F(256'hA0D6A9618580A9487FE961A5B2484C031002F0BC2B20F8177231800000008080),
       .INIT_50(256'hB86720B9A0E0A9E04320B9A0C1A9B85020B9A0BCA9BB0F20B9A0DBA9B86720B9),
       .INIT_51(256'h2070A5298528852785268500A9BAB720BA8B4C03D0BA8C20B9A0E5A9BD7E2068),
       .INIT_52(256'h094AB9834C03D0BB8F4CBA5E2062A5BA592063A5BA592064A5BA592065A5BA59),
       .INIT_53(256'h66266626856A6526A527856B6527A528856C6528A529856D6529A5181990A880),
       .INIT_54(256'h6B8522B1886C8522B1886D8522B104A02384228560D6D04A9870662966286627),
       .INIT_55(256'h04906165181FF069A56061A5698522B1886A8580096EA56F8566456E8522B188),
       .INIT_56(256'h4CB8F74C68680530FF4966A56066856FA5B8FB4C03D06185806914102C181D30),
       .INIT_57(256'h0C20000000208460E7F061E6B877206F8600A2F2B002691810F0AABC0C20B97E),
       .INIT_58(256'hB720618561E53800A9BC1B2076F0BA8C20BB124CBBA2206F8600A2BAA0F9A9BC),
       .INIT_59(256'h0865C46DA404D064C46CA40AD063C46BA410D062C46AA401A9FCA2BAF061E6BA),
       .INIT_5A(256'h6DA5A8E210CE30E6B06A266B266C266D060EB02801A9341032F02995E809902A),
       .INIT_5B(256'h0A0ACED040A9BB4F4C986A8562E56AA56B8563E56BA56C8564E56CA56D8565E5),
       .INIT_5C(256'h4C658529A5648528A5638527A5628526A5A4374C14A2BB8F4C2870850A0A0A0A),
       .INIT_5D(256'h8862858009668522B188638522B188648522B188658522B104A023842285B8D7),
       .INIT_5E(256'h9165A504A023842286BC1B204AA449A604F000A057A22C5CA2607084618522B1),
       .INIT_5F(256'h66856EA5607084229161A588229162257F0966A588229163A588229164A58822),
       .INIT_60(256'h06FBF061A5607086F9D0CA689560B506A2BC1B20607086F9D0CA609568B505A2),
       .INIT_61(256'h00A96285BC2B206001A902B0FFA92A66A509F061A5B9384CF2D0B96F20F79070),
       .INIT_62(256'hA025842485606646B8D24C6685708561866485658500A92AFF4962A588A26385),
       .INIT_63(256'h12D063C524B1C819D062C5800924B121D061E4C230664524B1C4F0AAC824B100),
       .INIT_64(256'h384AF061A5BC314CFF49029066A528F065E524B170C57FA9C80BD064C524B1C8),
       .INIT_65(256'h802966A5A8606884B999200610F9C961A28AB94D206885FFA9AA09106624A0E9),
       .INIT_66(256'hA0A92A8049668466A57084BC9B2020B0A0C961A5606884B9B020628562056246),
       .INIT_67(256'h2DC90F90FB10CA5D940AA200A060A86585648563856285B8D24C078565A56185),
       .INIT_68(256'h0EF0ABC9179000732030D045C92EF02EC95B9000732005D02BC904F0678604D0),
       .INIT_69(256'h494C5EE53800A90E1060245C90007320606607D004F02BC908F0AAC90AF02DC9),
       .INIT_6A(256'h5EC6BAE22007F0F9D05EE6BAFE20091012F05E855DE5385EA5C3505F245F66BD),
       .INIT_6B(256'h2048BD0A4CBD7E2030E93868BAE2205DE602105F2448BFB44C60013067A5F9D0),
       .INIT_6C(256'hB97E4C1130602464A909900AC95EA5B86A4C61A66F8566456EA5BC3C2068BC0C),
       .INIT_6D(256'h6B6E9EFD276B6E9EFD1FBC3E9BBD304C5E8530E9387A7100A0180A5E65180A0A),
       .INIT_6E(256'hA901A0AB1E4CBDDF20BC49203890A26386628539A63AA5BDDA20A3A071A90028),
       .INIT_6F(256'h09B002F080E000A9BF044C03D061A630A9C87184668500FF992DA90210662420),
       .INIT_70(256'h1002F0BC5B20BDA0B3A912101EF0BC5B20BDA0B8A95D85F7A9BA2820BDA0BDA9),
       .INIT_71(256'h0BC909300A69185DA501A2BC9B20B84920DCD05DE6BAFE20EED05DC6BAE2200E),
       .INIT_72(256'h30A906F08A00FF99C82EA971A4131002F08A5D865E8502E93802A9AAFF6906B0),
       .INIT_73(256'h6385BF177963A56485BF187964A56585BF19791865A580A200A0718400FF99C8),
       .INIT_74(256'hA44784C8C8C8C82F690A69FF4904908ADA300230DE1004B0E86285BF167962A5),
       .INIT_75(256'h04F024C0AA8029FF498A47A4718400FF99C82EA906D05DC600FF997F29AAC871),
       .INIT_76(256'h5EE53800A908102EF05EA62BA9C801F02EC9F8F030C98800FFB971A4A6D03CC0),
       .INIT_77(256'h9900A90102998A0103993A69FBB00AE9E8382FA28A01009945A90101992DA9AA),
       .INIT_78(256'hF0FF80969800001F0AFA00000000806001A000A901009900A900FF9908F00104),
       .INIT_79(256'h0300800ADFFFFFFFFFFF0A0000009CFFFFFFE8030000F0D8FFFFA0860100C0BD),
       .INIT_7A(256'hAAAAAAAAAAAAAAAAAAAAAAAAAAEC3C000000A8FDFFFF100E00006073FFFFC04B),
       .INIT_7B(256'hD069A570F0BBA220BFA011A9BC0C20AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA),
       .INIT_7C(256'hFE2007A49803D0BC5B2000A04EA9BCCC200F106EA5BBD42000A04EA2B8F94C03),
       .INIT_7D(256'h81606685FF4966A506F061A50A904A68BFED20BA282000A04EA9B9EA204898BB),
       .INIT_7E(256'h757E0A5859637C2A1C841D7A85E3EE2F771BB37E1674563E58347107293BAA38),
       .INIT_7F(256'hE0004CBC23200390506970A5BA2820BFA0BFA900000000811018723180C6E7FD),
       
       // The next set of INITP_xx are for the parity bits
       .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
       
       // The next set of INIT_xx are valid when configured as 36Kb
       .INITP_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0F(256'h0000000000000000000000000000000000000000000000000000000000000000)
    ) BRAM_SINGLE_MACRO_inst_BLOCK_1 (
       .DO(DATA_OUT_BLOCK_1),       // Output data, width defined by READ_WIDTH parameter
       .ADDR(addr[11:0]),   // Input address, width defined by read/write port depth
       .CLK(clk_counter[24]),     // 1-bit input clock
       .DI(0),       // Input data port, width defined by WRITE_WIDTH parameter
       .EN(1),       // 1-bit input RAM enable
       .REGCE(0), // 1-bit input output register enable
       .RST(0),     // 1-bit input reset
       .WE(8'h00)        // Input write enable, width defined by write port depth
    );
 
 
 //===============================================================================================
 
    BRAM_SINGLE_MACRO #(
       .BRAM_SIZE("36Kb"), // Target BRAM, "18Kb" or "36Kb" 
       .DEVICE("7SERIES"), // Target Device: "7SERIES" 
       .DO_REG(0), // Optional output register (0 or 1)
       .INIT(36'h000000000), // Initial values on output port
       .INIT_FILE ("NONE"),
       .WRITE_WIDTH(8), // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
       .READ_WIDTH(8),  // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
       .SRVAL(36'h000000000), // Set/Reset value for port output
       .WRITE_MODE("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE" 
       .INIT_00(256'h69B505A24801E938F3F081691807A5BCCC20BAD420039088C961A5BC0F205685),
       .INIT_01(256'h20686F8500A9E05920BFA0C4A9BFB420B85320708556A5F510CA6994619561B4),
       .INIT_02(256'hBBC72072847185BA284C00A057A9E05D20BA282057A9BBCA207284718560BAB9),
       .INIT_03(256'h847185C8019005691872A471A5BA282072A4718572E602D098C871A4678571B1),
       .INIT_04(256'hF32020D03730BC2B200046B12868007A44359860E4D067C600A05CA9B8672072),
       .INIT_05(256'h8BA9E0E34C658522B1C8638522B108A0648522B1C8628522B104A023842286FF),
       .INIT_06(256'h8564A563A66286658562A565A6B86720E0A092A9BA2820E0A08DA9BBA22000A0),
       .INIT_07(256'h86388407D0F0C9BBD44C00A08BA2B8D720618580A9708561A5668500A9648663),
       .INIT_08(256'hC62060DCB0E4AD2060E2B0FFCF2060E8B0FFD220A4374C1EA202D0AAA6634C37),
       .INIT_09(256'h030DAE030CAD48030FAD4846A948E1A9B7F720AD8A2060D0B0FFE42060D6B0FF),
       .INIT_0A(256'h202BA92EA42DA6E1D42060030F8D68030E8C030D8E030C8D0800146C28030EAC),
       .INIT_0B(256'h1CA217F00AA557B0FFD5202CA42BA60AA5E1D4200A8500A92C01A96095B0FFD8),
       .INIT_0C(256'h374C1DA205F0BF29FFB72060AB1E4CA3A064A907F002C97AA517D01029FFB720),
       .INIT_0D(256'h1920A6774CA53320A68E20A52A4CAB1E20A3A076A92E842D860ED002C97BA5A4),
       .INIT_0E(256'hFFBA2000A001A2FFBD2000A9E0F94CC390FFC32049A5E21920600BB0FFC020E2),
       .INIT_0F(256'hFFBA4C49A6A88AE20020E20620FFBA20498600A0E20020E20620E25720E20620),
       .INIT_10(256'h1120FFBD2000A9AF084CF7D0007920AEFD2060686802D0007920B79E4CE20E20),
       .INIT_11(256'h2088019003E049A500A04A86E20020E20620FFBA2000A001A28A4986B79E20E2),
       .INIT_12(256'hA422A6B6A320AD9E20E20E20E20620FFBA2049A54AA6A88AE20020E20620FFBA),
       .INIT_13(256'h8500A9BCCC20BC0C20BB07206EA6E2A0E5A9BC0C20B86720E2A0E0A9FFBD4C23),
       .INIT_14(256'hBFB4201285FF4912A5093066A5B849200D104866A5B85020E2A0EAA9B853206F),
       .INIT_15(256'h4EA2E26B20128500A9BBCA20E0434CE2A0EFA9BFB420031068B86720E2A0EAA9),
       .INIT_16(256'hE29D4C48BB0F4C00A04EA9E2DC2012A5668500A9BBA22000A057A9E0F62000A0),
       .INIT_17(256'h870189689987F8FB0728861B2D1AE68405000000007FA2DA0F4983A2DA0F4981),
       .INIT_18(256'hA0BCA9079081C94861A5BFB42003104866A5A2DA0F498328E75DA586E1DF3523),
       .INIT_19(256'h760B60BFB44C031068B85020E2A0E0A9079081C968E04320E3A03EA9BB0F20B9),
       .INIT_1A(256'hEAB77D4C7064147DC1CB53DE7CCA671F0C7C10B0FC837BF5A6F41E79D3BD83B3),
       .INIT_1B(256'h00A9FFCC20000000008113AAAAAA7FC791CC4C7E3A9944927E7E8830637D7A51),
       .INIT_1C(256'h9AFBA2E42220E3BF20E45320A4744CA43A4C03308A03006C80A258A67A201385),
       .INIT_1D(256'hA95852C74F8060D0E93830E938EFF020C90AB03AC9EA60AD7BE602D07AE6E4D0),
       .INIT_1E(256'h04840385B1A0AAA906840585B3A091A903128C03118DB2A048A903108D54854C),
       .INIT_1F(256'h19A201FC8E01FD8E01A218851385688500A9538503A9F810CA7395E3A2BD1CA2),
       .INIT_20(256'hE602D02BE62B919800A03484338638843786FF9920382C842B86FF9C20381686),
       .INIT_21(256'hA060A9BDCD202CE538A5AA2BE53837A5AB1E20E4A073A9A408202CA42BA5602C),
       .INIT_22(256'h0060F710CA03009DE447BD0BA2AE86A7E4A71AA57CA483E38BA6444CAB1E20E4),
       .INIT_23(256'h4F43202A2A2A2A202020200D93000D4545524620534554594220434953414220),
       .INIT_24(256'h52204B3436200D0D2A2A2A2A2032562043495341422034362045524F444F4D4D),
       .INIT_25(256'hAAAAAAAAAAAAAAAAAA608A019068AAFFC92048810020204D4554535953204D41),
       .INIT_26(256'h60F3910286AD60AB8501A9A985AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA),
       .INIT_27(256'h006900AE013702D106060C700DE8111A1944261960F7D0A1C504D0C891A40269),
       .INIT_28(256'h02918D00A9E5A02060D3A4D6A6E56C20D384D68607B06019A028A260DCA000A2),
       .INIT_29(256'h0CA9028B8D04A902868D0EA9028C8D02898D0AA902908DEBA9028F8D48A9CF85),
       .INIT_2A(256'h18A2D995FFA9F3D01AE0E8C80190286918D994AA00A9A880090288ADCC85CD85),
       .INIT_2B(256'hA9E9F020F410CAD3852869180830D9B4D3A5D6A6D684D38400A0FA10CAE9FF20),
       .INIT_2C(256'hE5664CE5A020EA60E6ED4C03F0C9E4EA244CD585F610E82869180630D9B4E827),
       .INIT_2D(256'hE802779D0278BD00A20277AC60F7D0CACFFF9DECB8BD2FA2998500A99A8503A9),
       .INIT_2E(256'h0287AECEA50CF0CFA578F7F002928DCC85C6A5E7162060185898C6C6F5D0C6E4),
       .INIT_2F(256'h0DC9CFF0F7D0CA02769DECE6BDC6867809A210D083C9E5B420EA1320CF8400A0),
       .INIT_30(256'hA61B30C9A5D484D38402928C00A0C884C8F7D08803D020C9D1B1D084D5A4C8D0),
       .INIT_31(256'hD785D1B1D3A493F0D0A5488A48982BB00A90C8C5D385CAA512D0C9E4E59120D6),
       .INIT_32(256'h8500A917D0C8C4E68420D3E64009027004D0D4A6049080090210D724D7063F29),
       .INIT_33(256'h02D0DEC9D7A5A868AA68D7850DA9E7162003F003E09AA606F003E099A60DA9D0),
       .INIT_34(256'hAED8C602F0D8A6800902F0C7A640096022A9D4850149D4A508D022C96018FFA9),
       .INIT_35(256'hB0D3C5D5A5D3E6E8B32060581868AA68D44602F0D8A5A868E6B620EA13200286),
       .INIT_36(256'hB5E8D956D916D6A6D6C6E8EA20079019E0D6A6E9674C03F00292AD32F04FC93F),
       .INIT_37(256'hD38500A9E87C20D6C6E9F04CF9D0CA0330D9B5D585286918D5A5CAD9958009D9),
       .INIT_38(256'h8500A94898488AD7854860D384D5A4E56C20D686CA9DD06868D38606D0D6A660),
       .INIT_39(256'h203F2902D0DF29049060C9109020C9E8914C03D00DC9E7D44C0310D7A5D3A4D0),
       .INIT_3A(256'h20D38488E8A120E7734CE7012006D0982ED014C9E6974C03F0D8A6E6934CE684),
       .INIT_3B(256'hD4A64D10F3910286ADD19120A9EFD0D5C4C8F39188F3B1C8D19188D1B1C8EA24),
       .INIT_3C(256'h90D5C488D384E8B320C817D01DC9E5662003D013C9C78502D012C9E6974C03F0),
       .INIT_3D(256'hD6C6EAF0EC90D5C5D6E6A8286998181DD011C9E6A84CD38400A0E87C20D6C609),
       .INIT_3E(256'h039020C95EA902D07FC97F29EC444CE8CB20E6A84CE87C20F8D0D385049028E9),
       .INIT_3F(256'h4FC007D0D3C404D020C9D1B1D5A437D014C93FD0D4A6E8914C03D00DC9E6914C),
       .INIT_40(256'hADD19120A9EFD0D3C488F391C8F3B188D191C8D1B188EA2420D5A4E9652024F0),
       .INIT_41(256'hE938D3A5D6C637F0D6A616D011C9E6974C400905F0D8A6E6A84CD8E6F3910286),
       .INIT_42(256'h8488E8A12009F09812D01DC9C78500A904D012C925D0E56C202A10D385049028),
       .INIT_43(256'hD6A6C946EC4F4CE8CB208009E6A84CE5442006D013C9E6A84CE70120E6A84CD3),
       .INIT_44(256'hA84CE87C20D386D486C786D88600A2E56C4CD686F410D9B5E8EA2003D019E0E8),
       .INIT_45(256'hD0CA28691807F0D3C527A902A260D6C660F6D0CA28691807F0D3C500A902A2E6),
       .INIT_46(256'h1E9C9F1C05906002868E60F810CA04F0E8DADD0FA260D6E602F019E0D6A660F6),
       .INIT_47(256'hE802A5CEC9C6D6C6FFA248AFA548AEA548ADA548ACA59B9A9998979695819E1F),
       .INIT_48(256'h0210DAB47F29D9B500A2E9FF20EC30E9C820DAB5AC85ECF1BD0CB018E0E9F020),
       .INIT_49(256'hDC01ADDC008D7FA902A5EED6E6C310D9A5F1858009F1A5EFD018E0E8D9958009),
       .INIT_4A(256'h8568AE8568AF8568D6A6C684F9D088FCD0CAEA00A00BD028DC008D7FA908FBC9),
       .INIT_4B(256'hDA4CD6C6CA02A5AEE8EA200C900EF018E002A58EFB10D9B5E8D6A660AC8568AD),
       .INIT_4C(256'hB5AC85ECEFBD0CF00E9002A5ECE9F020CA19A248AFA548AEA548ADA548ACA5E6),
       .INIT_4D(256'hAEECD0CADA9580090210D9B47F29DAB50F9002A5EC17A2E9FF20E930E9C820D8),
       .INIT_4E(256'h60F51088F391AEB1D191ACB127A0E9E020AD8502880D0329E9584CE6DA2002A5),
       .INIT_4F(256'hA060D28502880D0329D9B5D185ECF0BD60AF85D8090329ADA5AE85ACA5EA2420),
       .INIT_50(256'hD191D3A498EA2420CD8502A9A8EA60F61088D19120A9E4DA20EA2420E9F02027),
       .INIT_51(256'hCD8514A925D0CDC629D0CCA5FFEA2060F485D8090329D2A5F385D1A560F3918A),
       .INIT_52(256'h1C208049CEA50286AE02878DF3B1EA2420CE85CFE611B0D1B10287AECF46D3A4),
       .INIT_53(256'h0DADEA872001851F2901A506D0C0A508D0200901A5C08400A00AF0102901A5EA),
       .INIT_54(256'hA9F58581A9A861F0FFE0DC01AEDC008DCB8440A0028D8D00A94068AA68A868DC),
       .INIT_55(256'hF003C90CB005C9F5B14816B04AF8D0DC01CDDC01AD4808A2DC008DFEA9F685EB),
       .INIT_56(256'h028F6C68CCD0DC008D2A6838DFD0CA0BB041C0C868CB840210028D8D028D0D08),
       .INIT_57(256'hF014C929F07FC949701630028A2C7F2936D0028C8C10A007F0C5C4AAF5B1CBA4),
       .INIT_58(256'h8B8C04A026D0028BCE2BD0028CCE05F0028CAC35D011C904F01DC908F020C90C),
       .INIT_59(256'hE802779D06B00289ECC6A68A0EF0FFE0028E8C028DACC584CBA41C1088C6A402),
       .INIT_5A(256'h188D0249D018AD1D300291ADEEF0028ECD15D003C9028DAD60DC008D7FA9C686),
       .INIT_5B(256'h78EC03EBC2EB81EAE04CF685EB7ABDF585EB79BDAA06A9029008C90AEB764CD0),
       .INIT_5C(256'h5548423847593758544643364452350145535A3441573311878685881D0D14EC),
       .INIT_5D(256'h51022032045F312F5E3D01133B2A5C2C403A2E2D4C502B4E4F4B4D304A493956),
       .INIT_5E(256'hC8C228C7D927D8D4C6C326C4D22501C5D3DA24C1D723918B8A898C9D8D94FF03),
       .INIT_5F(256'h02A022045F213FDE3D01935DC0A93CBA5B3EDDCCD0DBCECFCBCD30CAC929D6D5),
       .INIT_60(256'hBF9BA5B79ABDA3BBBC99ACB29801B1AEAD97B0B396918B8A898C9D8D94FF83D1),
       .INIT_61(256'hA095045F813FDE3D01935DDFA83CA45B3EDCB6AFA6AAB9A1A730B5A229BEB8B4),
       .INIT_62(256'h08C9E6A84CD0188DFD29D018AD0BD08EC909D00209D018AD07D00EC9FF83AB02),
       .INIT_63(256'hFFFFFFFFFFFFFFFFE6A84C02918D02912D7FA9EED009C9093002910D80A907D0),
       .INIT_64(256'h0E0F0B0D920A0912161508029E07191F181406031E04129CFF05131A9F01171C),
       .INIT_65(256'h00000000000000FFFF11FFFF05FF0690FF1E1FFFFF1DFF1CFF001BFFFF0C10FF),
       .INIT_66(256'h0004030201060E0000000000000F140008000000379B00000000000000000000),
       .INIT_67(256'h583008E0B890684018F0C8A0785028000D4E55520D44414F4C07060504030201),
       .INIT_68(256'hA3469446ED4020A366380A10942448F0A42020092C4009C098704820F8D0A880),
       .INIT_69(256'hEEB320EE9720EE8E2078DD008D0809DD00ADEE852003D03FC9EE972078958568),
       .INIT_6A(256'h20FB90EEA920FBB0EEA920FB90EEA9200A10A324EE852064B0EEA920EE972078),
       .INIT_6B(256'hEE8520EE972003D0EEA02005B095663F900AF8D0DD00CDDD00ADA58508A9EE8E),
       .INIT_6C(256'hADDC0DADDC0F8D19A9DC078D04A9D4D0A5C6DD008D1009DF29DD00ADEAEAEAEA),
       .INIT_6D(256'h00ADED362095854A901858FE1C2003A92C80A96058F4B0EEA9200AD00229DC0D),
       .INIT_6E(256'h3094246058FB30EEA920EE8520EDBE20EEA02078ED3620958560DD008DF729DD),
       .INIT_6F(256'h3FA92C5FA9DD008D0809DD00ADEE8E20786018958568ED40204805D094663805),
       .INIT_70(256'hFB10EEA920EE8520A58500A978EE974CEE8520AAFDD0CA0AA28AEDBE20ED1120),
       .INIT_71(256'hA5A51810F430EEA92007D00229DC0DADDC0DADEE9720DC0F8D19A9DC078D01A9),
       .INIT_72(256'hDD00CDDD00ADA58508A9CAD0A5E6FE1C2040A9EE8520EEA020EDB24C02A905F0),
       .INIT_73(256'hEE062003509024EEA020E4D0A5C6F5300AF8D0DD00CDDD00ADA466F5100AF8D0),
       .INIT_74(256'h60DD008DDF29DD00AD60DD008D1009DD00AD60DD008DEF29DD00AD601858A4A5),
       .INIT_75(256'h3047F0B4A560AAFDD0CAB8A28A600AF8D0DD00CDDD00AD60DD008D2009DD00AD),
       .INIT_76(256'h1C3014F002942C20A960B58504298A06F0B4C6BD85BD458ACA019000A2B6463F),
       .INIT_77(256'hE650E970EAD0EDF0BDA5F0D0B4E6DFD0B4C6E3100293ADB4C6CA01D0BDA51470),
       .INIT_78(256'h9DACB4860298AEB585BD8500A91E501D10DD012C07904A0294ADCBD0FFA2B4E6),
       .INIT_79(256'hA14DDD0D8D01A902978D02970D10A92C40A960029DEEB685F9B113F0029ECC02),
       .INIT_7A(256'hF0A8C633D0A9A660CACA0250CA01F002932C20A909A260DD0D8D02A18D800902),
       .INIT_7B(256'h90A9EFD0A86501A90A0293AD67F0A7A5A8C660AA66A746AB85AB45A7A50D3036),
       .INIT_7C(256'h2AF0029CCCC8029BACE4D34CEAD0A7A5EF3B4C02A9A98502A18D02A10DDD0D8D),
       .INIT_7D(256'hAB45A7A5B130B4F002942C20A9F791F8D0E84A04F009E00298AEAAA588029B8C),
       .INIT_7E(256'hF0F1D0AAA5EF7E4C02978D02970D02A92C80A92C04A92C01A9A6502CA97003F0),
       .INIT_7F(256'h01ADFB70DD012CF9D0022902A1AD20D01D10DD012C02A929904A0294AD9A85EC),
       
       // The next set of INITP_xx are for the parity bits
       .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
       
       // The next set of INIT_xx are valid when configured as 36Kb
       .INITP_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0F(256'h0000000000000000000000000000000000000000000000000000000000000000)
    ) BRAM_SINGLE_MACRO_inst_BLOCK_2 (
       .DO(DATA_OUT_BLOCK_2),       // Output data, width defined by READ_WIDTH parameter
       .ADDR(addr[11:0]),   // Input address, width defined by read/write port depth
       .CLK(clk_counter[24]),     // 1-bit input clock
       .DI(0),       // Input data port, width defined by WRITE_WIDTH parameter
       .EN(1),       // 1-bit input RAM enable
       .REGCE(0), // 1-bit input output register enable
       .RST(0),     // 1-bit input reset
       .WE(8'h00)        // Input write enable, width defined by write port depth
    );
 
 
 //===============================================================================================
 
    BRAM_SINGLE_MACRO #(
       .BRAM_SIZE("36Kb"), // Target BRAM, "18Kb" or "36Kb" 
       .DEVICE("7SERIES"), // Target Device: "7SERIES" 
       .DO_REG(0), // Optional output register (0 or 1)
       .INIT(36'h000000000), // Initial values on output port
       .INIT_FILE ("NONE"),
       .WRITE_WIDTH(8), // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
       .READ_WIDTH(8),  // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
       .SRVAL(36'h000000000), // Set/Reset value for port output
       .WRITE_MODE("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE" 
       .INIT_00(256'hF4F0029DCCC8029EACF02820601802978D40A9F9300770DD012CDD018D0209DD),
       .INIT_01(256'hA9DD058D029AADDD048D0299ADDD0E8D10A91EB04A02A1ADF9919EA588029E8C),
       .INIT_02(256'hAD10DD012C02A924F0082928904A0294AD998560DD0E8D11A9EF0620EF3B2081),
       .INIT_03(256'h02A1ADEF3B4C1890A9F9F00429DD01ADDD018DFD29DD01ADFAB04A02A1AD22F0),
       .INIT_04(256'h978D080960029CEEF7B102978DF7290BF0029BCC029CAC0297AD6018F3F01229),
       .INIT_05(256'h2F490D606802A18D00A9DD0D8D10A9F9D0032902A1AD11F002A1AD486000A902),
       .INIT_06(256'h502053534552500DA0524F46A0474E494843524145530DA320524F525245204F),
       .INIT_07(256'h4F2059414C5020262044524F434552205353455250C5504154204E4F2059414C),
       .INIT_08(256'hC74E495946495245560DA0474E495641530DC74E4944414F4C0DC5504154204E),
       .INIT_09(256'h99A56018F31028C8FFD2207F2908F0BDB90D109D248D4B4F0DA0444E554F460D),
       .INIT_0A(256'hA5CA85D3A50BD099A5601897A4F08620978418D002C9E5B44C780FF0C6A508D0),
       .INIT_0B(256'h16B0F1992097863FF002C938B0E6324CC885D5A5D08509D003C9E6324CC985D6),
       .INIT_0C(256'h41200BD0F80D206097A68A68AA606897A6A6C6FE1C2040A905D00DB0F1992048),
       .INIT_0D(256'hD000C9F7B0F14E20EE134C60180DA904F090A56018B2B1F0F0A68500A911B0F8),
       .INIT_0E(256'h8A9E85684AEDDD4C680490E7164C6804D003C99AA548EEF0E9D060290297ADF2),
       .INIT_0F(256'h68A86818B2919EA5A684C8B29100A002A90EB0F864200ED0F80D202390489848),
       .INIT_10(256'hF003C916F0BAA5F31F20F7014C03F0F30F20F1FC4CF017206000A902909EA5AA),
       .INIT_11(256'h200610B9A5ED0920AA60189985F70A4C03F060E0B9A6F04D4C03D002C914B012),
       .INIT_12(256'h4C03D0BAA5F31F20F7014C03F0F30F20F7074CE61090248AEDC720F2484CEDCC),
       .INIT_13(256'h10B9A5ED0C20AA60189A85EAF060E0B9A6EFE14C03D002C911B00FF003C9F70D),
       .INIT_14(256'hF0BAA5488AF31F20601802F0F31420F7074CE71090248AEDB92003D0EDBE2005),
       .INIT_15(256'hA9C801F0FAA5C801F0F8A5FE2720F48320F2F220681DD002C947B04CF003C950),
       .INIT_16(256'h6000A9680490F86420F1DD203800A9F7D02023F00F29B9A5F47D4CFA85F88500),
       .INIT_17(256'h599D0259B998A414F098E498C6AA68F64220F2F14CF76A2005A90BD062C9B9A5),
       .INIT_18(256'hBD60F8D00259DD1530CA98A68A908500A96018026D9D026DB902639D0263B902),
       .INIT_19(256'h03B099E4EDFE2003B09AE403A2988500A960B985026DBDBA850263BDB8850259),
       .INIT_1A(256'h4C03900AE098A6F6FE4C03D0F30F20F70A4C03D0B8A660998500A99A86EDEF20),
       .INIT_1B(256'h20059056F003C95AF002639DBAA5026D9DB9856009B9A502599DB8A598E6F6FB),
       .INIT_1C(256'hAF2036B0F817201FD00F29B9A5F7134C03B0F7D020F4094C03D002C94F90F3D5),
       .INIT_1D(256'h2004A917B0F83820F4B00C9020F0F72C20F7044C28F01890F7EA200AF0B7A5F5),
       .INIT_1E(256'h8500A9F6F0B7A4FA30B9A56018A68598B29102A900A007F060C0B9A4BFA9F76A),
       .INIT_1F(256'hDD20BBB100A00CF0B7A5F7074C6868051090A5EDB920F009B9A5ED0C20BAA590),
       .INIT_20(256'hEF4A20F2D004C0C8029399BBB10AF0B7C402978CF48320F6544CF6D0B7C4C8ED),
       .INIT_21(256'hE4EABDE4EBBCF4404CFEC0BDFEC1BC09D002A6ADAA0A1CF00F290293AD02988E),
       .INIT_22(256'h8D029BADF00D2003B00ADD01AD09904A0294ADFF2E200A0295AD02958D02968C),
       .INIT_23(256'hF0A938F986FA848805D0FAA5F786F8848805D0F8A5FE2720029D8D029EAD029C),
       .INIT_24(256'hC3866002A18C00A0DD008DDD000D04A9DD018DDD038D06A9DD0D8D7FA9FE2D4C),
       .INIT_25(256'hA6F7104C03D0B7A47B90F9F003C9F7134C03D0BAA5908500A9938503306CC484),
       .INIT_26(256'h50B04A4A90A5AE85EE1320EDC720B9A5ED0920BAA5F3D520B98560A9F5AF20B9),
       .INIT_27(256'h334C03D0FFE12090859025FDA9F5D220AF85C4A5AE85C3A508D08AAF85EE1320),
       .INIT_28(256'hAEE6AE912CFE1C2010A908F0AED100A00CF093A48AE8B04A4A90A5AAEE1320F6),
       .INIT_29(256'h134C03B0F7D020F7134C03B04AF7044C7990F64220EDEF20CB509024AFE602D0),
       .INIT_2A(256'h2990A5D3B053F0F72C20DAB05AF00B90F7EA2009F0B7A5F5AF2068B0F81720F7),
       .INIT_2B(256'hB103A0EFD0B9A504B0C485B2B1C8C385B2B101A0DDD003E011F001E04AD03810),
       .INIT_2C(256'hC4A5C185C3A5AF85C46598AE85C3658A18A8B2F102A0B2B104A0AAB2F101A0B2),
       .INIT_2D(256'h2F2017A015F0B7A5F12F200CA01E109DA560AFA4AEA61824F84A20F5D220C285),
       .INIT_2E(256'h84AE86F12B4C59A002F093A549A060F6D0B7C4C8FFD220BBB100A00CF0B7A4F1),
       .INIT_2F(256'hB7A4B98561A95F90F9F003C9F7134C03D0BAA503326CC28501B5C18500B5AAAF),
       .INIT_30(256'hA5EDDD20ACA5FB8E2000A0EDB920B9A5ED0C20BAA5F68F20F3D520F7104C03D0),
       .INIT_31(256'h20E5D0FCDB20603800A9F6422007D0FFE120EDDD20ACB116B0FCD120EDDD20AD),
       .INIT_32(256'h20F7134C03B04A6018EDFE20EDB920E009EF29B9A5ED0C20BAA51130B924EDFE),
       .INIT_33(256'hB0F8672012B0F76A208A01A202D00129B9A503A2F68F2025B0F838208D90F7D0),
       .INIT_34(256'hD0A2E600A2F5C14CF12F2051A0FB109DA5601824F76A2005A906F00229B9A50D),
       .INIT_35(256'hCDDC01ADA286A186A08606904FE9A0A51AE9A1A501E9A2A538A0E602D0A1E606),
       .INIT_36(256'hA2A57860918502D0E8DC008DF8D0DC01ECDC01AEDC008EBDA21330AAF8D0DC01),
       .INIT_37(256'h02A92C01A96028C685FFCC200807D07FC991A56058A084A186A28578A0A4A1A6),
       .INIT_38(256'h200A509D2400A0FFCC204809A92C08A92C07A92C06A92C05A92C04A92C03A92C),
       .INIT_39(256'hC92AF005C9B2B100A032B0938568F841204893A5603868FFD22030094868F12F),
       .INIT_3A(256'hD015C0C8FFD220B2B105A0F12F2063A017109D24AAE1D004C904F003C908F001),
       .INIT_3B(256'hA9BFA048AEA548AFA548C1A548C2A55E90F7D0209E85608818EAE4E020A1A5F6),
       .INIT_3C(256'h84C8B291AFA5C8B291AEA5C8B291C2A5C8B291C1A5C8B2919EA5FBD088B29120),
       .INIT_3D(256'h6B20AB8569A9F7D720EED09FE69EE6B2919FA4BBB10CF0B7C49EA49E8400A09F),
       .INIT_3E(256'hC06918C1858AF7D0206002C0B3A4B2A66098C28568C18568AF8568AE8568A8F8),
       .INIT_3F(256'hD19FA4BBB110F0B7C49E8400A09F8405A01DB0F72C2060AF850069C28598AE85),
       .INIT_40(256'h2F201BA01AF0F82E2060C0C0A6A4A6E6F7D0206018ECD09EA49FE69EE6E7D0B2),
       .INIT_41(256'hD02EA0F9F0F82E206018012402D0012410A9F12F4C6AA0F8D0F82E20F8D020F1),
       .INIT_42(256'h90A99C859F859E85B085B485AA8500A9781FB0F81720F7D7209385908500A9DD),
       .INIT_43(256'hDC0EADDC0D8DDC0D8C7FA008A282A9786CB0F83820AB8514A9F7D72011D00EA2),
       .INIT_44(256'hA08D0315AD029F8D0314ADD0118DEF29D011ADF0A42002A28D9129DC0F8D1909),
       .INIT_45(256'hA0AD58F8D0CAFDD088FFA0FFA2C08501851F2901A5FB9720BE8502A9FCBD2002),
       .INIT_46(256'hA08D00A9686838FC93200BD018FFE120F8BE4CF6BC20F8D02015F0180315CD02),
       .INIT_47(256'h06ADAA2AB1062AB1062A0130B02400A9B185B16518B065180A0AB0A5B1866002),
       .INIT_48(256'hF01029DC0DAD02A48DDC0E8D02A2ADDC058DDC076D8ADC048DB165F99016C9DC),
       .INIT_49(256'hDC068CAAB186F2D0DC07ECDC06ED98FFA0DC07AE6058FF434C482AA948F9A909),
       .INIT_4A(256'hB1C53C6918B0A5B1664AB1664AB186B1E59802A38DDC0DADDC0F8D19A9DC078C),
       .INIT_4B(256'h17B0B1C5B0652669E81CB0B1C5B065306900A21B30A3A6FA604C03F09CA64AB0),
       .INIT_4C(256'h9265B1E513E938A9C602B0A9E619D0A8851DF0B4A5FA104C0390B1C5B0652C69),
       .INIT_4D(256'hA48500A916D002A4AD05D0012902A3AD22F0B4A5D7862BF0A4850149A4A59285),
       .INIT_4E(256'hB0E62CB0C6033007F092A5FEBC4CB9D09BA5F8E220A6A2BF303010A3A502A48D),
       .INIT_4F(256'hD2F0B4A59B859B458AB5B09685B99010C9BD30A9A5A0D08A0FD0D7E4928500A9),
       .INIT_50(256'h46F9974C0330A3A507F0B4A504F096A5FEBC4CF8E220DAA2BF66D746C530A3C6),
       .INIT_51(256'h8D81A9968500A9A88526F096A511D0B4A59CE6F8E220AA0AB065B1E53893A9B1),
       .INIT_52(256'hFEBC4CB685A905A8A5BD85BFA5DC0D8D01A9B48500A909F0B58596A5B485DC0D),
       .INIT_53(256'hA90BD0CABEA60CD0B5A51710AA240FA9A78502F0BEA5F8E220DAA29C85FB9720),
       .INIT_54(256'h0330BDA54AA7A5F1D0B6A5F5D0B5A518D03170FEBC4CAA8500A904D0FE1C2008),
       .INIT_55(256'hCAD0AA8580A9D0F0AB8500A9FB8E20AA8540A9DDD0AAC6AA850F2915B0181890),
       .INIT_56(256'hA00CF093A52DF0CAA7A6FB484C0390FCD120FB4A4C00A9FE1C2004A90AF0B5A5),
       .INIT_57(256'h009DACA501019DADA59EA63E909EE43DA24BF0B6A5B68501A904F0ACD1BDA500),
       .INIT_58(256'h9FE69FE627D00101DDADA52ED00100DDACA535F09EE49FA6FB3A4C9E86E8E801),
       .INIT_59(256'hA5A805D093A509D0FE1C2010A907F0B6A5B684C817F0ACD100A0BDA50BF093A5),
       .INIT_5A(256'h08F0A7C6BE860230CABEA6DC0DAEDC0D8E01A278AA8580A943D0FCDB20AC91BD),
       .INIT_5B(256'hF290FCD120FCDB20AB85AB45ACB1AB8400A0FB8E20FC932023F0BE8527D09EA5),
       .INIT_5C(256'h85A48500A9A38508A960AC85C1A5AD85C2A5FEBC4CFE1C2020A905F0BD45ABA5),
       .INIT_5D(256'hA5DC0F8D19A9DC0DADDC078EDC068D00A2B0A9029060A94ABDA560A9859B85A8),
       .INIT_5E(256'h2910B6A5A8E62FD0FBB12001A210A912D0A8A53C30B666386008290185084901),
       .INIT_5F(256'h49BDA50FF0A4850149A4A514D0FBA62019D0A9E61DD0FBAD2009D0A9A5FC574C),
       .INIT_60(256'h00A212F0A5A558FB9720F3103AF0A3A5A3C6BD46FEBC4C9B859B450129BD8501),
       .INIT_61(256'hA0CAB0BD85D7A5ADE691D00A90FCD120D9D0BD85800902D002E0BEA6A5C6D786),
       .INIT_62(256'h50A9FCCA2003D0BEC6FEBC4CBD8501499BA5BBD0FCDB20D785D745BD85ACB100),
       .INIT_63(256'hBD200AA2D810ABC6FB9720DFD0A7C6E3D0FBAF2078A9EAD0FCBD207808A2A785),
       .INIT_64(256'hFCCA20D0118D1009D011AD780883D0B686A58609A2FB8E2030F0BEA5ABE658FC),
       .INIT_65(256'hFD93BD97F0FC9320602803148D029FAD03158D09F002A0ADFDDD20DC0D8D7FA9),
       .INIT_66(256'hE602D0ACE660AFE5ADA5AEE5ACA538600185200901A56003158DFD94BD03148D),
       .INIT_67(256'h6C58FF5B20FD1520FD5020FDA320D0168E80006C03D0FD0220D89A78FFA260AD),
       .INIT_68(256'h1FA0C484C38618FDA030A23038CDC2C360F5D0CA03D08003DDFD0FBD05A2A000),
       .INIT_69(256'hF333F250F20EF291F34AFE47FE66EA3160F11088031499C391C3B102B00314B9),
       .INIT_6A(256'hA2F4D0C8030099020099000299A800A9F5EDF4A5FE66F32FF13EF6EDF1CAF157),
       .INIT_6B(256'h08D0C1D1C1912A0FD0C1D1C19155A9AAC1B1C2E6C28503A9A8B384B28603A03C),
       .INIT_6C(256'h31FBCDFC6A6002888D04A902828D08A9FE2D2018C2A4AA98E4F0E8D0C8C1918A),
       .INIT_6D(256'h038E00A2DD0F8DDC0F8DDD0E8DDC0E8D08A9DC008DDD0D8DDC0D8D7FA9F92CEA),
       .INIT_6E(256'h02A6AD00852FA90185E7A9DD028D3FA9DD008D07A9DC028ECAD4188EDD038EDC),
       .INIT_6F(256'h60BC84BB86B785FF6E4CDC058D42A9DC048D95A9FDF34C40A9DC048D25A90AF0),
       .INIT_70(256'h9085900590A59D85606802978D00A9480297AD0DD002C9BAA560B984BA86B885),
       .INIT_71(256'h8C02818E0282AC0281AE06906002848C02838E0284AC0283AE06906002858D60),
       .INIT_72(256'hBC2080026C03D0FD02201C30DD0DACDD0D8D7FA94898488A4803186C78600282),
       .INIT_73(256'hFB29DD00AD28F00129AA02A12D98A0026CE51820FDA320FD15200CD0FFE120F6),
       .INIT_74(256'hEEBB20FF0720FE9D4CFED62006F002290DF012298ADD0D8D02A1ADDD008DB505),
       .INIT_75(256'hAA68A868DD0D8D02A1ADFF072003F010298AFEB64CFED62006F002298AFEB64C),
       .INIT_76(256'hDD06ADA7850129DD01AD007100B8014602F006450CED0E7411C51A3E27C14068),
       .INIT_77(256'h068DFFA9DD0D8D02A1ADDD0F8D11A9DD078D029A6DDD07ADDD068D02996D1CE9),
       .INIT_78(256'h02A18D02A14D12A9DD0F8D11A9DD078D0296ADDD068D0295ADEF594CDD078DDD),
       .INIT_79(256'h029A8D00699802998DC8698AA82A0296ADAA60A8860298AEDD078DDD068DFFA9),
       .INIT_7A(256'h12ADE5182003146C03166C03F010290104BDBA4898488A4848EF296808EAEA60),
       .INIT_7B(256'hEE8E4CDC0E8D11098029DC0EADDC0D8D81A9FDDD4C02A68D0129D019ADFBD0D0),
       .INIT_7C(256'h4CFE344CFE254CEDC74CEDB94CFE184CFD1A4CFD154CFD504CFDA34CFF5B4C03),
       .INIT_7D(256'hFDF94CFE004CFE074CED094CED0C4CEDFE4CEDEF4CEDDD4CEE134CFE214CEA87),
       .INIT_7E(256'hDD4CF6E44CF5DD4CF49E4C03266C03246C03226C03206C031E6C031C6C031A6C),
       .INIT_7F(256'hFF48FCE2FE4359425252E5004CE50A4CE5054CF69B4C032C6C032A6C03286CF6),
       
       // The next set of INITP_xx are for the parity bits
       .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
       
       // The next set of INIT_xx are valid when configured as 36Kb
       .INITP_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0F(256'h0000000000000000000000000000000000000000000000000000000000000000)
    ) BRAM_SINGLE_MACRO_inst_BLOCK_3 (
       .DO(DATA_OUT_BLOCK_3),       // Output data, width defined by READ_WIDTH parameter
       .ADDR(addr[11:0]),   // Input address, width defined by read/write port depth
       .CLK(clk_counter[24]),     // 1-bit input clock
       .DI(0),       // Input data port, width defined by WRITE_WIDTH parameter
       .EN(1),       // 1-bit input RAM enable
       .REGCE(0), // 1-bit input output register enable
       .RST(0),     // 1-bit input reset
       .WE(8'h00)        // Input write enable, width defined by write port depth
    );
 
 
 //===============================================================================================
 
    BRAM_SINGLE_MACRO #(
       .BRAM_SIZE("36Kb"), // Target BRAM, "18Kb" or "36Kb" 
       .DEVICE("7SERIES"), // Target Device: "7SERIES" 
       .DO_REG(0), // Optional output register (0 or 1)
       .INIT(36'h000000000), // Initial values on output port
       .INIT_FILE ("NONE"),
       .WRITE_WIDTH(8), // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
       .READ_WIDTH(8),  // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
       .SRVAL(36'h000000000), // Set/Reset value for port output
       .WRITE_MODE("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE" 
       .INIT_00(256'h003C66606060663C007C66667C66667C006666667E663C18003C62606E6E663C),
       .INIT_01(256'h003C66666E60663C006060607860607E007E60607860607E00786C6666666C78),
       .INIT_02(256'h00666C7870786C6600386C0C0C0C0C1E003C18181818183C006666667E666666),
       .INIT_03(256'h003C66666666663C0066666E7E7E7666006363636B7F7763007E606060606060),
       .INIT_04(256'h003C66063C60663C00666C787C66667C000E3C666666663C006060607C66667C),
       .INIT_05(256'h0063777F6B63636300183C6666666666003C666666666666001818181818187E),
       .INIT_06(256'h003C30303030303C007E6030180C067E001818183C6666660066663C183C6666),
       .INIT_07(256'h0010307F7F301000181818187E3C1800003C0C0C0C0C0C3C00FC62307C30120C),
       .INIT_08(256'h006666FF66FF6666000000000066666600180000181818180000000000000000),
       .INIT_09(256'h0000000000180C06003F6667383C663C00466630180C666200187C063C603E18),
       .INIT_0A(256'h000018187E1818000000663CFF3C66000030180C0C0C1830000C18303030180C),
       .INIT_0B(256'h006030180C0603000018180000000000000000007E0000003018180000000000),
       .INIT_0C(256'h003C66061C06663C007E60300C06663C007E181818381818003C6666766E663C),
       .INIT_0D(256'h00181818180C667E003C66667C60663C003C6606067C607E0006067F661E0E06),
       .INIT_0E(256'h30181800001800000000180000180000003C66063E66663C003C66663C66663C),
       .INIT_0F(256'h001800180C06663C0070180C060C18700000007E007E0000000E18306030180E),
       .INIT_10(256'h000000FFFF0000001818181818181818003E1C7F7F3E1C08000000FFFF000000),
       .INIT_11(256'h30303030303030300000FFFF000000000000000000FFFF0000000000FFFF0000),
       .INIT_12(256'h000000E0F0381818000000070F1C1818181838F0E00000000C0C0C0C0C0C0C0C),
       .INIT_13(256'hC0C0C0C0C0C0FFFFC0E070381C0E070303070E1C3870E0C0FFFFC0C0C0C0C0C0),
       .INIT_14(256'h00081C3E7F7F7F3600FFFF0000000000003C7E7E7E7E3C00030303030303FFFF),
       .INIT_15(256'h003C7E66667E3C00C3E77E3C3C7EE7C318181C0F070000006060606060606060),
       .INIT_16(256'h181818FFFF18181800081C3E7F3E1C080606060606060606003C181866661818),
       .INIT_17(256'h0103070F1F3F7FFF003636763E03000018181818181818183030C0C03030C0C0),
       .INIT_18(256'h00000000000000FFFFFFFFFF00000000F0F0F0F0F0F0F0F00000000000000000),
       .INIT_19(256'h03030303030303033333CCCC3333CCCCC0C0C0C0C0C0C0C0FF00000000000000),
       .INIT_1A(256'h1818181F1F181818030303030303030380C0E0F0F8FCFEFF3333CCCC00000000),
       .INIT_1B(256'hFFFF000000000000181818F8F80000000000001F1F1818180F0F0F0F00000000),
       .INIT_1C(256'h181818F8F8181818181818FFFF000000000000FFFF1818181818181F1F000000),
       .INIT_1D(256'h000000000000FFFF0707070707070707E0E0E0E0E0E0E0E0C0C0C0C0C0C0C0C0),
       .INIT_1E(256'hF0F0F0F000000000FFFF030303030303FFFFFF00000000000000000000FFFFFF),
       .INIT_1F(256'h0F0F0F0FF0F0F0F000000000F0F0F0F0000000F8F8181818000000000F0F0F0F),
       .INIT_20(256'hFFC3999F9F9F99C3FF83999983999983FF9999998199C3E7FFC3999F919199C3),
       .INIT_21(256'hFFC39999919F99C3FF9F9F9F879F9F81FF819F9F879F9F81FF87939999999387),
       .INIT_22(256'hFF9993878F879399FFC793F3F3F3F3E1FFC3E7E7E7E7E7C3FF99999981999999),
       .INIT_23(256'hFFC39999999999C3FF99999181818999FF9C9C9C9480889CFF819F9F9F9F9F9F),
       .INIT_24(256'hFFC399F9C39F99C3FF99938783999983FFF1C399999999C3FF9F9F9F83999983),
       .INIT_25(256'hFF9C8880949C9C9CFFE7C39999999999FFC3999999999999FFE7E7E7E7E7E781),
       .INIT_26(256'hFFC3CFCFCFCFCFC3FF819FCFE7F3F981FFE7E7E7C3999999FF9999C3E7C39999),
       .INIT_27(256'hFFEFCF8080CFEFFFE7E7E7E781C3E7FFFFC3F3F3F3F3F3C3FF039DCF83CFEDF3),
       .INIT_28(256'hFF99990099009999FFFFFFFFFF999999FFE7FFFFE7E7E7E7FFFFFFFFFFFFFFFF),
       .INIT_29(256'hFFFFFFFFFFE7F3F9FFC09998C7C399C3FFB999CFE7F3999DFFE783F9C39FC1E7),
       .INIT_2A(256'hFFFFE7E781E7E7FFFFFF99C300C399FFFFCFE7F3F3F3E7CFFFF3E7CFCFCFE7F3),
       .INIT_2B(256'hFF9FCFE7F3F9FCFFFFE7E7FFFFFFFFFFFFFFFFFF81FFFFFFCFE7E7FFFFFFFFFF),
       .INIT_2C(256'hFFC399F9E3F999C3FF819FCFF3F999C3FF81E7E7E7C7E7E7FFC39999899199C3),
       .INIT_2D(256'hFFE7E7E7E7F39981FFC39999839F99C3FFC399F9F9839F81FFF9F98099E1F1F9),
       .INIT_2E(256'hCFE7E7FFFFE7FFFFFFFFE7FFFFE7FFFFFFC399F9C19999C3FFC39999C39999C3),
       .INIT_2F(256'hFFE7FFE7F3F999C3FF8FE7F3F9F3E78FFFFFFF81FF81FFFFFFF1E7CF9FCFE7F1),
       .INIT_30(256'hFFFFFF0000FFFFFFE7E7E7E7E7E7E7E7FFC1E38080C1E3F7FFFFFF0000FFFFFF),
       .INIT_31(256'hCFCFCFCFCFCFCFCFFFFF0000FFFFFFFFFFFFFFFFFF0000FFFFFFFFFF0000FFFF),
       .INIT_32(256'hFFFFFF1F0FC7E7E7FFFFFFF8F0E3E7E7E7E7C70F1FFFFFFFF3F3F3F3F3F3F3F3),
       .INIT_33(256'h3F3F3F3F3F3F00003F1F8FC7E3F1F8FCFCF8F1E3C78F1F3F00003F3F3F3F3F3F),
       .INIT_34(256'hFFF7E3C1808080C9FF0000FFFFFFFFFFFFC381818181C3FFFCFCFCFCFCFC0000),
       .INIT_35(256'hFFC381999981C3FF3C1881C3C381183CE7E7E3F0F8FFFFFF9F9F9F9F9F9F9F9F),
       .INIT_36(256'hE7E7E70000E7E7E7FFF7E3C180C1E3F7F9F9F9F9F9F9F9F9FFC3E7E79999E7E7),
       .INIT_37(256'hFEFCF8F0E0C08000FFC9C989C1FCFFFFE7E7E7E7E7E7E7E7CFCF3F3FCFCF3F3F),
       .INIT_38(256'hFFFFFFFFFFFFFF0000000000FFFFFFFF0F0F0F0F0F0F0F0FFFFFFFFFFFFFFFFF),
       .INIT_39(256'hFCFCFCFCFCFCFCFCCCCC3333CCCC33333F3F3F3F3F3F3F3F00FFFFFFFFFFFFFF),
       .INIT_3A(256'hE7E7E7E0E0E7E7E7FCFCFCFCFCFCFCFC7F3F1F0F07030100CCCC3333FFFFFFFF),
       .INIT_3B(256'h0000FFFFFFFFFFFFE7E7E70707FFFFFFFFFFFFE0E0E7E7E7F0F0F0F0FFFFFFFF),
       .INIT_3C(256'hE7E7E70707E7E7E7E7E7E70000FFFFFFFFFFFF0000E7E7E7E7E7E7E0E0FFFFFF),
       .INIT_3D(256'hFFFFFFFFFFFF0000F8F8F8F8F8F8F8F81F1F1F1F1F1F1F1F3F3F3F3F3F3F3F3F),
       .INIT_3E(256'h0F0F0F0FFFFFFFFF0000FCFCFCFCFCFC000000FFFFFFFFFFFFFFFFFFFF000000),
       .INIT_3F(256'hF0F0F0F00F0F0F0FFFFFFFFF0F0F0F0FFFFFFF0707E7E7E7FFFFFFFFF0F0F0F0),
       .INIT_40(256'h003C6060603C0000007C66667C606000003E663E063C0000003C62606E6E663C),
       .INIT_41(256'h7C063E66663E0000001818183E180E00003C607E663C0000003E66663E060600),
       .INIT_42(256'h00666C786C6060003C06060606000600003C181838001800006666667C606000),
       .INIT_43(256'h003C6666663C000000666666667C000000636B7F7F660000003C181818183800),
       .INIT_44(256'h007C063C603E000000606060667C000006063E66663E000060607C66667C0000),
       .INIT_45(256'h00363E7F6B63000000183C6666660000003E666666660000000E1818187E1800),
       .INIT_46(256'h003C30303030303C007E30180C7E0000780C3E666666000000663C183C660000),
       .INIT_47(256'h0010307F7F301000181818187E3C1800003C0C0C0C0C0C3C00FC62307C30120C),
       .INIT_48(256'h006666FF66FF6666000000000066666600180000181818180000000000000000),
       .INIT_49(256'h0000000000180C06003F6667383C663C00466630180C666200187C063C603E18),
       .INIT_4A(256'h000018187E1818000000663CFF3C66000030180C0C0C1830000C18303030180C),
       .INIT_4B(256'h006030180C0603000018180000000000000000007E0000003018180000000000),
       .INIT_4C(256'h003C66061C06663C007E60300C06663C007E181818381818003C6666766E663C),
       .INIT_4D(256'h00181818180C667E003C66667C60663C003C6606067C607E0006067F661E0E06),
       .INIT_4E(256'h30181800001800000000180000180000003C66063E66663C003C66663C66663C),
       .INIT_4F(256'h001800180C06663C0070180C060C18700000007E007E0000000E18306030180E),
       .INIT_50(256'h003C66606060663C007C66667C66667C006666667E663C18000000FFFF000000),
       .INIT_51(256'h003C66666E60663C006060607860607E007E60607860607E00786C6666666C78),
       .INIT_52(256'h00666C7870786C6600386C0C0C0C0C1E003C18181818183C006666667E666666),
       .INIT_53(256'h003C66666666663C0066666E7E7E7666006363636B7F7763007E606060606060),
       .INIT_54(256'h003C66063C60663C00666C787C66667C000E3C666666663C006060607C66667C),
       .INIT_55(256'h0063777F6B63636300183C6666666666003C666666666666001818181818187E),
       .INIT_56(256'h181818FFFF181818007E6030180C067E001818183C6666660066663C183C6666),
       .INIT_57(256'h66CC993366CC9933CCCC3333CCCC333318181818181818183030C0C03030C0C0),
       .INIT_58(256'h00000000000000FFFFFFFFFF00000000F0F0F0F0F0F0F0F00000000000000000),
       .INIT_59(256'h03030303030303033333CCCC3333CCCCC0C0C0C0C0C0C0C0FF00000000000000),
       .INIT_5A(256'h1818181F1F1818180303030303030303663399CC663399CC3333CCCC00000000),
       .INIT_5B(256'hFFFF000000000000181818F8F80000000000001F1F1818180F0F0F0F00000000),
       .INIT_5C(256'h181818F8F8181818181818FFFF000000000000FFFF1818181818181F1F000000),
       .INIT_5D(256'h000000000000FFFF0707070707070707E0E0E0E0E0E0E0E0C0C0C0C0C0C0C0C0),
       .INIT_5E(256'hF0F0F0F000000000006070786C060301FFFFFF00000000000000000000FFFFFF),
       .INIT_5F(256'h0F0F0F0FF0F0F0F000000000F0F0F0F0000000F8F8181818000000000F0F0F0F),
       .INIT_60(256'hFFC39F9F9FC3FFFFFF839999839F9FFFFFC199C1F9C3FFFFFFC3999F919199C3),
       .INIT_61(256'h83F9C19999C1FFFFFFE7E7E7C1E7F1FFFFC39F8199C3FFFFFFC19999C1F9F9FF),
       .INIT_62(256'hFF999387939F9FFFC3F9F9F9F9FFF9FFFFC3E7E7C7FFE7FFFF999999839F9FFF),
       .INIT_63(256'hFFC3999999C3FFFFFF9999999983FFFFFF9C94808099FFFFFFC3E7E7E7E7C7FF),
       .INIT_64(256'hFF83F9C39FC1FFFFFF9F9F9F9983FFFFF9F9C19999C1FFFF9F9F83999983FFFF),
       .INIT_65(256'hFFC9C180949CFFFFFFE7C3999999FFFFFFC199999999FFFFFFF1E7E7E781E7FF),
       .INIT_66(256'hFFC3CFCFCFCFCFC3FF81CFE7F381FFFF87F3C1999999FFFFFF99C3E7C399FFFF),
       .INIT_67(256'hFFEFCF8080CFEFFFE7E7E7E781C3E7FFFFC3F3F3F3F3F3C3FF039DCF83CFEDF3),
       .INIT_68(256'hFF99990099009999FFFFFFFFFF999999FFE7FFFFE7E7E7E7FFFFFFFFFFFFFFFF),
       .INIT_69(256'hFFFFFFFFFFE7F3F9FFC09998C7C399C3FFB999CFE7F3999DFFE783F9C39FC1E7),
       .INIT_6A(256'hFFFFE7E781E7E7FFFFFF99C300C399FFFFCFE7F3F3F3E7CFFFF3E7CFCFCFE7F3),
       .INIT_6B(256'hFF9FCFE7F3F9FCFFFFE7E7FFFFFFFFFFFFFFFFFF81FFFFFFCFE7E7FFFFFFFFFF),
       .INIT_6C(256'hFFC399F9E3F999C3FF819FCFF3F999C3FF81E7E7E7C7E7E7FFC39999899199C3),
       .INIT_6D(256'hFFE7E7E7E7F39981FFC39999839F99C3FFC399F9F9839F81FFF9F98099E1F1F9),
       .INIT_6E(256'hCFE7E7FFFFE7FFFFFFFFE7FFFFE7FFFFFFC399F9C19999C3FFC39999C39999C3),
       .INIT_6F(256'hFFE7FFE7F3F999C3FF8FE7F3F9F3E78FFFFFFF81FF81FFFFFFF1E7CF9FCFE7F1),
       .INIT_70(256'hFFC3999F9F9F99C3FF83999983999983FF9999998199C3E7FFFFFF0000FFFFFF),
       .INIT_71(256'hFFC39999919F99C3FF9F9F9F879F9F81FF819F9F879F9F81FF87939999999387),
       .INIT_72(256'hFF9993878F879399FFC793F3F3F3F3E1FFC3E7E7E7E7E7C3FF99999981999999),
       .INIT_73(256'hFFC39999999999C3FF99999181818999FF9C9C9C9480889CFF819F9F9F9F9F9F),
       .INIT_74(256'hFFC399F9C39F99C3FF99938783999983FFF1C399999999C3FF9F9F9F83999983),
       .INIT_75(256'hFF9C8880949C9C9CFFE7C39999999999FFC3999999999999FFE7E7E7E7E7E781),
       .INIT_76(256'hE7E7E70000E7E7E7FF819FCFE7F3F981FFE7E7E7C3999999FF9999C3E7C39999),
       .INIT_77(256'h993366CC993366CC3333CCCC3333CCCCE7E7E7E7E7E7E7E7CFCF3F3FCFCF3F3F),
       .INIT_78(256'hFFFFFFFFFFFFFF0000000000FFFFFFFF0F0F0F0F0F0F0F0FFFFFFFFFFFFFFFFF),
       .INIT_79(256'hFCFCFCFCFCFCFCFCCCCC3333CCCC33333F3F3F3F3F3F3F3F00FFFFFFFFFFFFFF),
       .INIT_7A(256'hE7E7E7E0E0E7E7E7FCFCFCFCFCFCFCFC99CC663399CC6633CCCC3333FFFFFFFF),
       .INIT_7B(256'h0000FFFFFFFFFFFFE7E7E70707FFFFFFFFFFFFE0E0E7E7E7F0F0F0F0FFFFFFFF),
       .INIT_7C(256'hE7E7E70707E7E7E7E7E7E70000FFFFFFFFFFFF0000E7E7E7E7E7E7E0E0FFFFFF),
       .INIT_7D(256'hFFFFFFFFFFFF0000F8F8F8F8F8F8F8F81F1F1F1F1F1F1F1F3F3F3F3F3F3F3F3F),
       .INIT_7E(256'h0F0F0F0FFFFFFFFFFF9F8F8793F9FCFE000000FFFFFFFFFFFFFFFFFFFF000000),
       .INIT_7F(256'hF0F0F0F00F0F0F0FFFFFFFFF0F0F0F0FFFFFFF0707E7E7E7FFFFFFFFF0F0F0F0),
       
       // The next set of INITP_xx are for the parity bits
       .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
       
       // The next set of INIT_xx are valid when configured as 36Kb
       .INITP_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0F(256'h0000000000000000000000000000000000000000000000000000000000000000)
    ) BRAM_SINGLE_MACRO_inst_BLOCK_4 (
       .DO(DATA_OUT_BLOCK_4),       // Output data, width defined by READ_WIDTH parameter
       .ADDR(addr[11:0]),   // Input address, width defined by read/write port depth
       .CLK(clk_counter[24]),     // 1-bit input clock
       .DI(0),       // Input data port, width defined by WRITE_WIDTH parameter
       .EN(1),       // 1-bit input RAM enable
       .REGCE(0), // 1-bit input output register enable
       .RST(0),     // 1-bit input reset
       .WE(8'h00)        // Input write enable, width defined by write port depth
    );
 
 
 //===============================================================================================
    
//    always clk = #10 ~clk;
    
    always @(posedge clk_counter[24])
    //if (!reset)
    begin
      addr <= addr + 1;
    end
    
    always @*
    case (addr[14:12])
      3'b000: combined_data_out = DATA_OUT_BLOCK_0;
      3'b001: combined_data_out = DATA_OUT_BLOCK_1;
      3'b010: combined_data_out = DATA_OUT_BLOCK_2;         
      3'b011: combined_data_out = DATA_OUT_BLOCK_3;
      3'b100: combined_data_out = DATA_OUT_BLOCK_4;
      default:  combined_data_out = 0;
    endcase
    
    always @(posedge clk_out)
    clk_counter <= clk_counter + 1; 
    
    
endmodule
