`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05.07.2017 15:35:00
// Design Name: 
// Module Name: test
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module rom_basic(
  input clk,
  input [12:0] addr,
  output DO
    );
    
    
    
    wire [7:0] DATA_OUT_BLOCK_0;
    wire [7:0] DATA_OUT_BLOCK_1;
    wire nc_wire;
    reg [7:0] combined_data_out;
    reg bit_12_store;
 
   BRAM_SINGLE_MACRO #(
       .BRAM_SIZE("36Kb"), // Target BRAM, "18Kb" or "36Kb" 
       .DEVICE("7SERIES"), // Target Device: "7SERIES" 
       .DO_REG(0), // Optional output register (0 or 1)
       .INIT(36'h000000000), // Initial values on output port
       .INIT_FILE ("NONE"),
       .WRITE_WIDTH(8), // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
       .READ_WIDTH(8),  // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
       .SRVAL(36'h000000000), // Set/Reset value for port output
       .WRITE_MODE("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE" 
       .INIT_00(256'hA89FA9A4AC05B080ABBEABA4A8F7AD1DA741A83043495341424D4243E37BE394),
       .INIT_01(256'hAA9FAA7FB823B3B2E164E155E167B82CA94AA82EA93AA8D1A882A81CA927A870),
       .INIT_02(256'hBF71B39EB37D0310BC58BCCCBC39A641AB7AE1C6E1BDE129AA85A65DA69BA856),
       .INIT_03(256'hB737B72CB700B6ECB78BB7ADB465B77CB80DE30EE2B4E26BE264BFEDB9EAE097),
       .INIT_04(256'h4E45B01564AED35ABFB37DAFE546AFE850BF7A7FBB117BBA2A7BB85279B86979),
       .INIT_05(256'h454CC4414552CD4944D455504E49A35455504E49C1544144D458454ED24F46C4),
       .INIT_06(256'h53CD4552CE5255544552C255534F47C5524F54534552C649CE5552CF544F47D4),
       .INIT_07(256'h5250C54B4F50C64544D94649524556C5564153C4414F4CD4494157CE4FD04F54),
       .INIT_08(256'h4C43CE45504FD35953C44D43D24C43D453494CD44E4F43D44E495250A3544E49),
       .INIT_09(256'hD0455453D44F4ECE454854A8435053CE46CF54A8424154D7454ED44547C5534F),
       .INIT_0A(256'h53D34F50C55246D25355D34241D44E49CE4753BCBDBED24FC44E41DEAFAAADAB),
       .INIT_0B(256'h5453CE454CCB454550CE5441CE4154CE4953D34F43D05845C74F4CC44E52D251),
       .INIT_0C(256'h4F5400CF47A444494DA45448474952A45446454CA4524843C35341CC4156A452),
       .INIT_0D(256'h504F20544F4E20454C4946CE45504F20454C4946D3454C494620594E414D204F),
       .INIT_0E(256'h455345525020544F4E20454349564544C44E554F4620544F4E20454C4946CE45),
       .INIT_0F(256'h4DC54C49462054555054554F20544F4EC54C4946205455504E4920544F4ED44E),
       .INIT_10(256'h4E20454349564544204C4147454C4C49C54D414E20454C494620474E49535349),
       .INIT_11(256'h5255544552D841544E5953D24F462054554F48544957205458454ED245424D55),
       .INIT_12(256'h4147454C4C49C154414420464F2054554FC255534F472054554F48544957204E),
       .INIT_13(256'h55D9524F4D454D20464F2054554FD74F4C465245564FD95449544E415551204C),
       .INIT_14(256'h444552D4504952435342555320444142D44E454D45544154532044274645444E),
       .INIT_15(256'h4147454C4C49CF52455A205942204E4F495349564944D9415252412044274D49),
       .INIT_16(256'h204F4F5420474E49525453C84354414D53494D2045505954D44345524944204C),
       .INIT_17(256'hD8454C504D4F43204F4F5420414C554D524F46C154414420454C4946C74E4F4C),
       .INIT_18(256'h4556CE4F4954434E55462044274645444E55C5554E49544E4F432054274E4143),
       .INIT_19(256'hA23BA235A225A210A1FFA1F0A1E2A1D0A1C2A1B5A1ACA19EC4414F4CD9464952),
       .INIT_1A(256'hA31EA30EA300A2EDA2E4A2D5A2C8A2BAA2AAA29DA290A27FA272A26AA25AA24F),
       .INIT_1B(256'h0A0D2E59444145520A0D00204E492000524F5252452020000D4B4F0DA383A324),
       .INIT_1C(256'hBD49850102BD0AD04AA521D081C90101BDE8E8E8E8BAA0004B414552420A0D00),
       .INIT_1D(256'h3832843185A4082060D8D0AA1269188A07F00102DD49A507D00103DD4A850103),
       .INIT_1E(256'h22E558A5385BC603B05A8522E5385AA523F098E8AA60E55BA5A822855FE55AA5),
       .INIT_1F(256'h35B03E690A60F2D0CA59C65BC658915AB1F9D08858915AB1049059C608B05885),
       .INIT_20(256'hA2B52620FA10CA57B5489809A248229033C504D0289034C4602E9022E4BA2285),
       .INIT_21(256'hA326BDAA0A8A03006C10A26001B033C505D0069034C468A868FA30E8619568F7),
       .INIT_22(256'h68C8AB47207F294822B100A0AB4520AAD720138500A9FFCC202385A327BD2285),
       .INIT_23(256'hFF902080A9AB1E20A3A076A9BDC22003F0C83AA4AB1E20A3A069A9A67A20F410),
       .INIT_24(256'h20A96B20A7E14CA5792006903A86FFA2F0F0AA0073207B847A86A5602003026C),
       .INIT_25(256'h852D65185FF1885FA5258560A522852DA523855FB101A04490A613200B84A579),
       .INIT_26(256'hB11823C6039022651825C6E803B0A82DE55FA538AA60E52E85FF692EA524852D),
       .INIT_27(256'h850B655A852DA51888F00200ADA53320A65920F2D0CA25E623E6F9D0C8249122),
       .INIT_28(256'hA42E842D8532A431A501FF8C01FE8D15A414A5A3B8205984C801905B842EA458),
       .INIT_29(256'h22B101A018238422852CA42BA5A4804CA53320A65920F810885F9101FCB9880B),
       .INIT_2A(256'h60DD90238522862291C8006923A5229100A0AA226598C8FBD022B1C804A01DF0),
       .INIT_2B(256'h04A07AA603046CAACA4CA4374C17A2F19059E0E802009D0DF00DC9E1122000A2),
       .INIT_2C(256'h04D03FC92D700F2456F022C9088537F020C9F4D0E83EF0FFC907100200BD0F84),
       .INIT_2D(256'hF0A09EF9380200BDE8C8CA7A86880B8400A071841D903CC9049030C925D099A9),
       .INIT_2E(256'hE9380F8502D049C904F03AE93836F001FBB901FB99C8E871A40B0530D080C9F5),
       .INIT_2F(256'hB9FA10A09DB9C80BE67AA6F0D0E801FB99C8DBF008C5DFF00200BD08859FD055),
       .INIT_30(256'hF05FB160865F8501A02CA62BA5607A85FFA97BC601FD99BE100200BDB4D0A09E),
       .INIT_31(256'hD7B05FB188AA5FB1880AF00C905FD18814A509D08803F018905FD115A5C8C81F),
       .INIT_32(256'h2DD000A9A68E202E8500692CA52D850269182BA52B91C82B91A800A9FDD06018),
       .INIT_33(256'hA868168619A2A81D203284318530842F852EA42DA53484338538A437A5FFE720),
       .INIT_34(256'h04F00690607B85FF692CA57A85FF692BA5186010853E8500A94898489AFAA268),
       .INIT_35(256'h0514A5686886D0A96B200073208ED0ABC90CF0007920A61320A96B20E9D0ABC9),
       .INIT_36(256'h15C55FB1C8AA5FB1C8AAD720A82C2043F05FB10F8401A015851485FFA906D015),
       .INIT_37(256'h0F85FF490FA506D022C9AB47207F2949A420A9BDCD2049842CB002F014E404D0),
       .INIT_38(256'hD3F0FFC9D71003066CE3864CB5D060855F865FB1C8AA5FB1A810D05FB111F0C8),
       .INIT_39(256'hAB4720B230A09EB9C8F530FA10A09EB9C808F0CAFFA04984AA7FE938CF300F24),
       .INIT_3A(256'h659818A90620A3FB2009A968689AAA0F698A05D0A38A20A9A520108580A9F5D0),
       .INIT_3B(256'h628562257F0966A5AD8A20AD8D20AEFF20A4A94839A5483AA54800697BA5487A),
       .INIT_3C(256'h20AD8A2000732006D0A9C9007920BBA220B9A0BCA9AE434C23842285A7A08BA9),
       .INIT_3D(256'h00A03E843D8504F0EA02C07BA47AA5A82C204881A94849A5484AA5AE3820BC2B),
       .INIT_3E(256'hE602907A857A65983A857AB1C839857AB1C8A84B4C03D0187AB102A043D07AB1),
       .INIT_3F(256'hA00CB948A00DB9A80A17B023C9119080E93CF0A7AE4CA7ED2000732003086C7B),
       .INIT_40(256'h2BA538A8A04CAEFF20A4A9007320F9D04BC9AF084CD6F03AC9A9A54C00734C48),
       .INIT_41(256'h843D850CF0E83AA67BA47AA53CD01801B0FFE12060428441858801B02CA401E9),
       .INIT_42(256'h4C03D03EA41AA217D0E3864CA4694C0390A3A081A968683C843B853AA439A53E),
       .INIT_43(256'hA66020A6594C03D028FF902000A908603A8439853CA43BA57B847A853DA5A437),
       .INIT_44(256'hA7AE4CA8A020007920488DA94839A5483AA5487AA5487BA5A3FB2003A9A8974C),
       .INIT_45(256'h2CA62BA504B0E807907BA67A6538980BB015E53AA514E539A538A90920A96B20),
       .INIT_46(256'h0BF08DC99AA38A204A85FFA9FDD0607B8500E960A57A8501E95FA51E90A61720),
       .INIT_47(256'h857A651898A906207B85687A85683A856839856868AF084CA4374C11A22C0CA2),
       .INIT_48(256'hF008C5E8F07AB10886078507A608A5088400A0078600A22C3AA2607BE602907A),
       .INIT_49(256'hBBF0A9092005D061A5AEFF20A7A905F089C9007920AD9E20E9F0F3D022C9C8E4),
       .INIT_4A(256'h20A7EF4C6804D065C691D089C904F08DC948B79E20A7ED4CA8A04C03B0007920),
       .INIT_4B(256'hA5D4B019C9228515A507852FE9F7B01586148600A26068EEF02CC9A96B200073),
       .INIT_4C(256'h2015E602901485076514A5152614061585156522A51485146522260A22260A14),
       .INIT_4D(256'hD0AD90202A68AD9E20480DA5480EA5AEFF20B2A94A844985B08B20A9714C0073),
       .INIT_4E(256'h4CD0BFC04AA468BBD04C60499165A5C8499164A500A0B1BF20BC1B2012106818),
       .INIT_4F(256'hAABC0C20AA1D2071A471E6BAE220AA1D2071846684618400A03DD006C9B6A620),
       .INIT_50(256'h2022B1FFDB4C65A563A464A6BC9B20BAE220DFD006C0C871A4BAED208AE805F0),
       .INIT_51(256'hC465A40E9033C564B18807D0179034C564B102A0BD7E4C2FE9B2484C03900080),
       .INIT_52(256'h846F8551A450A5B4752064B100A0AA684C65A464A507B02DC564A50DD008902E),
       .INIT_53(256'h60499150B1C8499150B1C8499150B100A0B6DB205184508500A061A9B67A2070),
       .INIT_54(256'h007920AB2120AAA04C28E11820138608AEFF202CA905F0B79E20ABB54CAA8620),
       .INIT_55(256'h20BDDD20DE300D24AD9E205EF03BC937F02CC94BF018A6C950F0A3C943F035F0),
       .INIT_56(256'h05101324AB47200DA910D013A501A0FFA202009D00A9D3D0AB3B20AB2120B487),
       .INIT_57(256'h200984FFF020380816D00169FF49FCB00AE93898FFF0203860FF49AB47200AA9),
       .INIT_58(256'h8720F2D0AB3B20AAA24C00732006D0CAE8AA059009E58A06902859D029C9B79B),
       .INIT_59(256'hA903F013A5AB284CAAE520F3D00DC9C8AB472022B1BCF0CAE800A0AAB6A620B4),
       .INIT_5A(256'h4C3A84398540A43FA504D0FFA0043011F011A560FF29E10C203FA92C1DA92C20),
       .INIT_5B(256'h23C9B3A620607B847A853EA43DA5AB1E20ADA00CA9A4374C18A205F013A5AF08),
       .INIT_5C(256'hAC0F2040A902018D00A902A001A2E11E201386AEFF202CA9B79E2000732010D0),
       .INIT_5D(256'hC960138600A2FFCC2013A5ABCE20E11E201386AEFF202CA9B79E206013D013A6),
       .INIT_5E(256'hFFB7200DF013A5ABF92001FF8D2CA9B3A620AB2120AEFF203BA9AEBD200BD022),
       .INIT_5F(256'hAB452006D013A5A8FB4CA90620E3D013A51ED00200ADA8F84CABB52006F00229),
       .INIT_60(256'h7BA47AA54A844985B08B2044844386118500A92C98A942A441A6A5604CAB3B20),
       .INIT_61(256'hD001A0FFA202008DE124200C50112420D00079207B847A8644A443A64C844B85),
       .INIT_62(256'hA97A86E80950112431100D240073207B847A86ABF920AB452003D013A575300C),
       .INIT_63(256'hB48D20C8019000697BA47AA50885182CA907853AA907F022C907850CF0078500),
       .INIT_64(256'hA47AA5AB4D4C03F02CC907F0007920A9C2200EA5BCF320AC914CA9DA20B7E220),
       .INIT_65(256'hA212D0AAC8A90620AC154CAEFD202DF00079207B847A854CA44BA5448443857B),
       .INIT_66(256'hA5AC514CDCD083E0AA007920A8FB204085C87AB1C83F857AB1C86CF07AB1C80D),
       .INIT_67(256'h5458453F60AB1E4CACA0FCA907D013A50BF043B100A0A8274C031011A644A443),
       .INIT_68(256'h04D0000D5452415453204D4F5246204F4445523F000D4445524F4E4749204152),
       .INIT_69(256'h6824850669480469188A9AA4374C0AA205F0A38A204A844985B08B2003F000A0),
       .INIT_6A(256'hF00109FD38BABC5D2001A0BBD020B867204AA449A566850109BDBABBA22001A0),
       .INIT_6B(256'h0079209AAA11698AA7AE4C7B850111BD7A850112BD3A850110BD3985010FBD17),
       .INIT_6C(256'h7AA6A4374C16A2FDB06003B003300D24382418AD9E20AD2420007320F1D02CC9),
       .INIT_6D(256'h1790B1E9380079204D8500A9AE8320A3FB2001A9488A482400A27AC67BC602D0),
       .INIT_6E(256'h9007697BB02CD04DA6ADBB4C0073204D8561904DC54D4501492A01C913B003C9),
       .INIT_6F(256'h4BA468AE202048AD8D2067B0A080D968A822650A2285FF69B63D4C03D00D6577),
       .INIT_70(256'hD99048B0A080D9D7D04D851BA07AC67BC602D07AA62A8A0D465FD056F0AA1710),
       .INIT_71(256'h856822E6228568A8A080BE66A5AF084CADA94C4DA5AE332048A081B948A082B9),
       .INIT_72(256'hF064C923F068FFA000226C4861A54862A54863A54864A54865A5BC1B20489823),
       .INIT_73(256'h6F8566456E85686D85686C85686B85686A856869856812854A684B84AD8D2003),
       .INIT_74(256'hA8A90FD0FFC9AF284C0390B11320BCF34C03B00073200D8500A9030A6C6061A5),
       .INIT_75(256'hA47AA50FD022C9D1F0AAC958F0ABC9DEF02EC9A1DA0F498200734CBBA220AEA0),
       .INIT_76(256'hFF4964A5A8FF4965A5B1BF203BD018A013D0A8C9B7E24CB48720C8019000697B),
       .INIT_77(256'hA02CA92C28A92C29A9AD9E20AEFA20AFA74C0390B4C9B3F44C03D0A5C9B3914C),
       .INIT_78(256'hA90890A0E965A500E964A538ADFA4C686815A0A4374C0BA200734C03D07AD100),
       .INIT_79(256'h1C90AF1420708500A926F00DA546A445A665846485B08B206065E5E3A964E5A2),
       .INIT_7A(256'h100E2460B46F4CBE682024A05D8406A07184885E84AF842014D0C9C018D054E0),
       .INIT_7B(256'hA298AF842025D049C01BD054E02D90AF1420B3914C8AA864B1C8AA64B100A00D),
       .INIT_7C(256'hBC3C4CFFB72006D054C00AD053E060628400A0658563846486FFDE20BC4F4CA0),
       .INIT_7D(256'hA5AA68AD8F20AEFD20AD9E20AEFA2020908FE0007320AA480ABBA24C65A464A5),
       .INIT_7E(256'h56859FEBB955859FEAB9A868AEF120AFD64C488AA868B79E20488A4864A54865),
       .INIT_7F(256'h20BBFC2008850B4565A507850B4564A5B1BF200B8400A02CFFA0AD8D4C005420),
       
       // The next set of INITP_xx are for the parity bits
       .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
       
       // The next set of INIT_xx are valid when configured as 36Kb
       .INITP_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0F(256'h0000000000000000000000000000000000000000000000000000000000000000)
    ) BRAM_SINGLE_MACRO_inst_BLOCK_0 (
       .DO(DATA_OUT_BLOCK_0),       // Output data, width defined by READ_WIDTH parameter
       .ADDR(addr[11:0]),   // Input address, width defined by read/write port depth
       .CLK(clk),     // 1-bit input clock
       .DI(0),       // Input data port, width defined by WRITE_WIDTH parameter
       .EN(1),       // 1-bit input RAM enable
       .REGCE(0), // 1-bit input output register enable
       .RST(0),     // 1-bit input reset
       .WE(8'h00)        // Input write enable, width defined by write port depth
    );
 
 
 //===============================================================================================
 
    BRAM_SINGLE_MACRO #(
       .BRAM_SIZE("36Kb"), // Target BRAM, "18Kb" or "36Kb" 
       .DEVICE("7SERIES"), // Target Device: "7SERIES" 
       .DO_REG(0), // Optional output register (0 or 1)
       .INIT(36'h000000000), // Initial values on output port
       .INIT_FILE ("NONE"),
       .WRITE_WIDTH(8), // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
       .READ_WIDTH(8),  // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
       .SRVAL(36'h000000000), // Set/Reset value for port output
       .WRITE_MODE("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE" 
       .INIT_00(256'h257F096EA513B0AD9020B3914C0B4507250B4564A5A80B4508250B4565A5B1BF),
       .INIT_01(256'hA46CA5638462866185B6A6204DC60D8500A9B0614CAABC5B2000A069A96A856A),
       .INIT_02(256'hA607D0CAC8E8FFA06685FFA961A6049001A908F061E538AA6D846C86B6AA206D),
       .INIT_03(256'hFD20BC3C4CFFA902F012252A8AE801A202B0FFA2EFF062D16CB10C90180F3066),
       .INIT_04(256'hA2AF084C03B0B1132000792045850C8600792000A260F4D0007920B09020AAAE),
       .INIT_05(256'hFFA906D024C9F6B0B11320FB90007320AA0B90B1132005900073200E860D8600),
       .INIT_06(256'h1005384686007320AA80098A458545050E8580A9D0D010A513D025C910D00D85),
       .INIT_07(256'hD05FD145A522F02FC504D030E45F8560862EA62DA5108400A0B1D14C03D028E9),
       .INIT_08(256'hC9486860A5E9385BE9059041C9DCD0E8E19007695FA518887DF05FD1C846A508),
       .INIT_09(256'hC004D053C9AF084C03D049C0EFF0C9C00BD054C946A445A560BFA013A905D02A),
       .INIT_0A(256'hA3B82059845885C801900769185B845A8532A431A560845F8530A42FA5F5F054),
       .INIT_0B(256'hC85F91C85F91C85F91C800A95F9146A5C85F9145A500A030842F85C859A458A5),
       .INIT_0C(256'hC8019060A45F6505690A0BA56048844785C8019060A40269185FA55F91C85F91),
       .INIT_0D(256'hA50D3066A5AD8D20AD9E200073206065A464A5B1BF2000000080906059845885),
       .INIT_0E(256'h4846A5489800A0480DA5480E050CA5BC9B4C7AD0BC5B20B1A0A5A9099090C961),
       .INIT_0F(256'h019D65A501029D64A5480101BD480102BDBAA868468568458568B1B2204845A5),
       .INIT_10(256'h60855F8630A52FA60C857F290E85680D8568AEF7200B84D2F02CC9007920C801),
       .INIT_11(256'hB1C8AA5F65185FB1C816F05FD146A506D045C5C85FB100A039F031E404D032C5),
       .INIT_12(256'hEA4CE7D05FD104A00BA5B19420F7D00CA513A2A4374C0EA22C12A2D79060655F),
       .INIT_13(256'hA57186CACA02105F9146A5C8CA01105F9145A505A2728400A0A40820B19420B2),
       .INIT_14(256'hB34C205F918AC85F91C8006968AA0169186808500C2400A90BA25F91C8C8C80B),
       .INIT_15(256'h32843185A4082052F0C8039058658AA859855DB05965DCD00BC622A472857186),
       .INIT_16(256'h32A55F9102A05FE531A53859E6F5D072C659C6FBD058918805F071A472E600A9),
       .INIT_17(256'h0E905FD16585686485AA68C87285718500A90B855FB1C862D00CA55F9160E5C8),
       .INIT_18(256'h22A498AA64658AB34C200AF018710572A5C8A4354CB2454C07905FD18AC806D0),
       .INIT_19(256'h658AB3552000A92886CACA021046A5CA011045A505A27285CAD00BC671866565),
       .INIT_1A(256'h8A00A000A25D8510A929855FB18828855FB122846047A5A84885596598478558),
       .INIT_1B(256'hF00DA560E3D05DC693B0A8296598AA28658A180B9072267106A4B0A82A98AA0A),
       .INIT_1C(256'h2038BC444C90A2638462850D8600A232E534A5A831E533A538B52620B6A62003),
       .INIT_1D(256'h108580A9AEFA20B3A620B3E120A4374C1BA22C15A2A0D0E83AA6EBF000A9FFF0),
       .INIT_1E(256'h4F4CA8F820487AA5487BA54847A54848A548AEFF20B2A9AEF720AD8D20B08B20),
       .INIT_1F(256'hAEF120484EA5484FA5B3E120AD8D4C4F844E85B0922010858009AEFF20A5A9B4),
       .INIT_20(256'h48A4FA10884847B1C8488599F04EB1C8AA47854EB102A04F85684E8568AD8D20),
       .INIT_21(256'h85684E8568AD8A204847A54848A57B854EB1C87A854EB1487AA5487BA5BBD420),
       .INIT_22(256'h4E91C8684E91C8684E91C8684E916800A07B85687A8568AF084C03F00079204F),
       .INIT_23(256'hB4F4205184508665A464A612F000A0FFA96868BDDF2000A0AD8D20604E91C868),
       .INIT_24(256'h04F007C50CF06FB1C8FFA06384628570846F850886078622A260618563846286),
       .INIT_25(256'h980BD002C904F070A57286E8019070A671856F659861841801F022C9F3D008C5),
       .INIT_26(256'h9563A5019562A5009561A5A4374C19A205D022E016A6B6882070A46FA6B47520),
       .INIT_27(256'h01B034A4336538FF49480F46601686E8E8E817860D848870846584648600A002),
       .INIT_28(256'hA9B52620B6300FA510A26068AA36843585348433850B9031C504D0119032C488),
       .INIT_29(256'h00A219A960865F8532A631A54E844F8400A03485338638A537A6D0D0680F8580),
       .INIT_2A(256'hF02FC504D030E4238622852EA62DA5538507A9F7F0B5C72005F016C523862285),
       .INIT_2B(256'h862285B6064C03D031C507D032E459A658A5538503A959865885F3F0B5BD2005),
       .INIT_2C(256'hB1C8D0308AD310285985596522B1C85885586522B1C80822B1C8AA22B100A023),
       .INIT_2D(256'h3022B1F3F0B5C720BAF058C504D059E423A623E602902285226505690A00A022),
       .INIT_2E(256'h169060C51AB033E41ED0069034C522B1C8AA22B1C82BF022B1C8301022B1C835),
       .INIT_2F(256'hE60290228522651853A5558553A54F864E8523A622A560855F8610905FE404D0),
       .INIT_30(256'h5B85006960A55A855F654EB15585A84A042955A5F5F04E054FA56000A023A623),
       .INIT_31(256'h4865A5B52A4C4E91C859A559E6AA4E9158A5C855A4A3BF205986588534A633A5),
       .INIT_32(256'hB47520A4374C17A205906471186FB100A07085686F8568AD8F20AE83204864A5),
       .INIT_33(256'hC8486FB100A0ADB84CB4CA20B6AA2070A46FA5B68C20B6AA2051A450A5B67A20),
       .INIT_34(256'h0290358535651868F8D098359122B188480AF0A82384228668A86FB1C8AA6FB1),
       .INIT_35(256'h68A822B1C8AA22B1C84822B100A008B6DB202384228565A464A5AD8F206036E6),
       .INIT_36(256'hC50CD018C460238422866834E602903385336518480BD033E40FD034C413D028),
       .INIT_37(256'hB4CA4C6868629100A068B47D2001A9488AB7A1206000A0178503E9168508D017),
       .INIT_38(256'h8522651868A868B6AA2051A450A5B47D20488A4898AA50B104909850D1B76120),
       .INIT_39(256'h29C90079206585FFA9B7064CFF4950F118B76120B4CA4CB68C209823E6029022),
       .INIT_3A(256'hB065A5B19065C5FF49B6B050F100A218488ACA4BF0B76120B79E20AEFD2006F0),
       .INIT_3B(256'h4CB78220608A00A048984855A5518568508568AA686868558568A868AEF720AD),
       .INIT_3C(256'h8A20007320B2484CB3A24CA822B100A008F0B7822060A80D8600A2B6A320B3A2),
       .INIT_3D(256'h8622A6728471867BA47AA6B8F74C03D0B7822000794C65A6F0D064A6B1B820AD),
       .INIT_3E(256'h00A068BCF3200079202491984824B100A02586E801907B8623A624852265187A),
       .INIT_3F(256'hB091C961A59D3066A5B79E4CAEFD20B7F720AD8A20607B847A8672A471A62491),
       .INIT_40(256'h8568148568A814B100A0B7F7204814A54815A5601585148465A464A5BC9B2097),
       .INIT_41(256'h00A04A86B7F12003F000792000A24986B7EB2060149100A08AB7EB20B3A24C15),
       .INIT_42(256'h4C61A56F856E456685FF4966A5BA8C20B8674CBFA011A960F8F049254A4514B1),
       .INIT_43(256'h9024F061E538CEF0A869A569A2568670A6BBFC4C03D0BA8C203C90B99920B86A),
       .INIT_44(256'h015670A5A8C730F9C9708400A004D061A2568400A00069FF4966846EA4618412),
       .INIT_45(256'h0003B9658504F50004B970855665FF493869A002F069E061A057106F24B9B020),
       .INIT_46(256'hA64AD062A6189800A0B9472003B0628501F50001B9638502F50002B9648503F5),
       .INIT_47(256'h5665606685618500A9E4D020C908697084658670A6648665A6638664A6628663),
       .INIT_48(256'h060169B9364C62856A6562A563856B6563A564856C6564A565856D6565A57085),
       .INIT_49(256'h6366626642F061E60E9061850169FF49C7B061E538F210622663266426652670),
       .INIT_4A(256'hA56485FF4964A56385FF4963A56285FF4962A56685FF4966A560706665666466),
       .INIT_4B(256'h0FA26062E602D063E606D064E60AD065E60ED070E67085FF4970A56585FF4965),
       .INIT_4C(256'hE9E6F0E8300869019468A4029401B4039402B4049403B4708404B425A2A4374C),
       .INIT_4D(256'h000000816018ECD0C86A0476037602760176017601F60290011614B070A5A808),
       .INIT_4E(256'h34F304358134F3043580203BAA38821693387680640B9B138079CB565E7F0300),
       .INIT_4F(256'hA0D6A9618580A9487FE961A5B2484C031002F0BC2B20F8177231800000008080),
       .INIT_50(256'hB86720B9A0E0A9E04320B9A0C1A9B85020B9A0BCA9BB0F20B9A0DBA9B86720B9),
       .INIT_51(256'h2070A5298528852785268500A9BAB720BA8B4C03D0BA8C20B9A0E5A9BD7E2068),
       .INIT_52(256'h094AB9834C03D0BB8F4CBA5E2062A5BA592063A5BA592064A5BA592065A5BA59),
       .INIT_53(256'h66266626856A6526A527856B6527A528856C6528A529856D6529A5181990A880),
       .INIT_54(256'h6B8522B1886C8522B1886D8522B104A02384228560D6D04A9870662966286627),
       .INIT_55(256'h04906165181FF069A56061A5698522B1886A8580096EA56F8566456E8522B188),
       .INIT_56(256'h4CB8F74C68680530FF4966A56066856FA5B8FB4C03D06185806914102C181D30),
       .INIT_57(256'h0C20000000208460E7F061E6B877206F8600A2F2B002691810F0AABC0C20B97E),
       .INIT_58(256'hB720618561E53800A9BC1B2076F0BA8C20BB124CBBA2206F8600A2BAA0F9A9BC),
       .INIT_59(256'h0865C46DA404D064C46CA40AD063C46BA410D062C46AA401A9FCA2BAF061E6BA),
       .INIT_5A(256'h6DA5A8E210CE30E6B06A266B266C266D060EB02801A9341032F02995E809902A),
       .INIT_5B(256'h0A0ACED040A9BB4F4C986A8562E56AA56B8563E56BA56C8564E56CA56D8565E5),
       .INIT_5C(256'h4C658529A5648528A5638527A5628526A5A4374C14A2BB8F4C2870850A0A0A0A),
       .INIT_5D(256'h8862858009668522B188638522B188648522B188658522B104A023842285B8D7),
       .INIT_5E(256'h9165A504A023842286BC1B204AA449A604F000A057A22C5CA2607084618522B1),
       .INIT_5F(256'h66856EA5607084229161A588229162257F0966A588229163A588229164A58822),
       .INIT_60(256'h06FBF061A5607086F9D0CA689560B506A2BC1B20607086F9D0CA609568B505A2),
       .INIT_61(256'h00A96285BC2B206001A902B0FFA92A66A509F061A5B9384CF2D0B96F20F79070),
       .INIT_62(256'hA025842485606646B8D24C6685708561866485658500A92AFF4962A588A26385),
       .INIT_63(256'h12D063C524B1C819D062C5800924B121D061E4C230664524B1C4F0AAC824B100),
       .INIT_64(256'h384AF061A5BC314CFF49029066A528F065E524B170C57FA9C80BD064C524B1C8),
       .INIT_65(256'h802966A5A8606884B999200610F9C961A28AB94D206885FFA9AA09106624A0E9),
       .INIT_66(256'hA0A92A8049668466A57084BC9B2020B0A0C961A5606884B9B020628562056246),
       .INIT_67(256'h2DC90F90FB10CA5D940AA200A060A86585648563856285B8D24C078565A56185),
       .INIT_68(256'h0EF0ABC9179000732030D045C92EF02EC95B9000732005D02BC904F0678604D0),
       .INIT_69(256'h494C5EE53800A90E1060245C90007320606607D004F02BC908F0AAC90AF02DC9),
       .INIT_6A(256'h5EC6BAE22007F0F9D05EE6BAFE20091012F05E855DE5385EA5C3505F245F66BD),
       .INIT_6B(256'h2048BD0A4CBD7E2030E93868BAE2205DE602105F2448BFB44C60013067A5F9D0),
       .INIT_6C(256'hB97E4C1130602464A909900AC95EA5B86A4C61A66F8566456EA5BC3C2068BC0C),
       .INIT_6D(256'h6B6E9EFD276B6E9EFD1FBC3E9BBD304C5E8530E9387A7100A0180A5E65180A0A),
       .INIT_6E(256'hA901A0AB1E4CBDDF20BC49203890A26386628539A63AA5BDDA20A3A071A90028),
       .INIT_6F(256'h09B002F080E000A9BF044C03D061A630A9C87184668500FF992DA90210662420),
       .INIT_70(256'h1002F0BC5B20BDA0B3A912101EF0BC5B20BDA0B8A95D85F7A9BA2820BDA0BDA9),
       .INIT_71(256'h0BC909300A69185DA501A2BC9B20B84920DCD05DE6BAFE20EED05DC6BAE2200E),
       .INIT_72(256'h30A906F08A00FF99C82EA971A4131002F08A5D865E8502E93802A9AAFF6906B0),
       .INIT_73(256'h6385BF177963A56485BF187964A56585BF19791865A580A200A0718400FF99C8),
       .INIT_74(256'hA44784C8C8C8C82F690A69FF4904908ADA300230DE1004B0E86285BF167962A5),
       .INIT_75(256'h04F024C0AA8029FF498A47A4718400FF99C82EA906D05DC600FF997F29AAC871),
       .INIT_76(256'h5EE53800A908102EF05EA62BA9C801F02EC9F8F030C98800FFB971A4A6D03CC0),
       .INIT_77(256'h9900A90102998A0103993A69FBB00AE9E8382FA28A01009945A90101992DA9AA),
       .INIT_78(256'hF0FF80969800001F0AFA00000000806001A000A901009900A900FF9908F00104),
       .INIT_79(256'h0300800ADFFFFFFFFFFF0A0000009CFFFFFFE8030000F0D8FFFFA0860100C0BD),
       .INIT_7A(256'hAAAAAAAAAAAAAAAAAAAAAAAAAAEC3C000000A8FDFFFF100E00006073FFFFC04B),
       .INIT_7B(256'hD069A570F0BBA220BFA011A9BC0C20AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA),
       .INIT_7C(256'hFE2007A49803D0BC5B2000A04EA9BCCC200F106EA5BBD42000A04EA2B8F94C03),
       .INIT_7D(256'h81606685FF4966A506F061A50A904A68BFED20BA282000A04EA9B9EA204898BB),
       .INIT_7E(256'h757E0A5859637C2A1C841D7A85E3EE2F771BB37E1674563E58347107293BAA38),
       .INIT_7F(256'hE0004CBC23200390506970A5BA2820BFA0BFA900000000811018723180C6E7FD),
       
       // The next set of INITP_xx are for the parity bits
       .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
       
       // The next set of INIT_xx are valid when configured as 36Kb
       .INITP_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
       .INITP_0F(256'h0000000000000000000000000000000000000000000000000000000000000000)
    ) BRAM_SINGLE_MACRO_inst_BLOCK_1 (
       .DO(DATA_OUT_BLOCK_1),       // Output data, width defined by READ_WIDTH parameter
       .ADDR(addr[11:0]),   // Input address, width defined by read/write port depth
       .CLK(clk),     // 1-bit input clock
       .DI(0),       // Input data port, width defined by WRITE_WIDTH parameter
       .EN(1),       // 1-bit input RAM enable
       .REGCE(0), // 1-bit input output register enable
       .RST(0),     // 1-bit input reset
       .WE(8'h00)        // Input write enable, width defined by write port depth
    );
 
 //===============================================================================================
    
    always @(posedge clk)
    bit_12_store <= addr[12];
       
    always @*
    case (bit_12_store)
      1'b0: combined_data_out = DATA_OUT_BLOCK_0;
      1'b1: combined_data_out = DATA_OUT_BLOCK_1;
      default:  combined_data_out = 0;
    endcase
   
    assign DO = combined_data_out;
    
endmodule
