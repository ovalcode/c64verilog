`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05.07.2017 15:35:00
// Design Name: 
// Module Name: test
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module rom_chargen(
  input clk,
  input [11:0] addr,
  output DO
  );
  
  
  
  wire [7:0] DATA_OUT_BLOCK_0;
  wire nc_wire;  

    BRAM_SINGLE_MACRO #(
     .BRAM_SIZE("36Kb"), // Target BRAM, "18Kb" or "36Kb" 
     .DEVICE("7SERIES"), // Target Device: "7SERIES" 
     .DO_REG(0), // Optional output register (0 or 1)
     .INIT(36'h000000000), // Initial values on output port
     .INIT_FILE ("NONE"),
     .WRITE_WIDTH(8), // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
     .READ_WIDTH(8),  // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
     .SRVAL(36'h000000000), // Set/Reset value for port output
     .WRITE_MODE("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE" 
     .INIT_00(256'h003C66606060663C007C66667C66667C006666667E663C18003C62606E6E663C),
     .INIT_01(256'h003C66666E60663C006060607860607E007E60607860607E00786C6666666C78),
     .INIT_02(256'h00666C7870786C6600386C0C0C0C0C1E003C18181818183C006666667E666666),
     .INIT_03(256'h003C66666666663C0066666E7E7E7666006363636B7F7763007E606060606060),
     .INIT_04(256'h003C66063C60663C00666C787C66667C000E3C666666663C006060607C66667C),
     .INIT_05(256'h0063777F6B63636300183C6666666666003C666666666666001818181818187E),
     .INIT_06(256'h003C30303030303C007E6030180C067E001818183C6666660066663C183C6666),
     .INIT_07(256'h0010307F7F301000181818187E3C1800003C0C0C0C0C0C3C00FC62307C30120C),
     .INIT_08(256'h006666FF66FF6666000000000066666600180000181818180000000000000000),
     .INIT_09(256'h0000000000180C06003F6667383C663C00466630180C666200187C063C603E18),
     .INIT_0A(256'h000018187E1818000000663CFF3C66000030180C0C0C1830000C18303030180C),
     .INIT_0B(256'h006030180C0603000018180000000000000000007E0000003018180000000000),
     .INIT_0C(256'h003C66061C06663C007E60300C06663C007E181818381818003C6666766E663C),
     .INIT_0D(256'h00181818180C667E003C66667C60663C003C6606067C607E0006067F661E0E06),
     .INIT_0E(256'h30181800001800000000180000180000003C66063E66663C003C66663C66663C),
     .INIT_0F(256'h001800180C06663C0070180C060C18700000007E007E0000000E18306030180E),
     .INIT_10(256'h000000FFFF0000001818181818181818003E1C7F7F3E1C08000000FFFF000000),
     .INIT_11(256'h30303030303030300000FFFF000000000000000000FFFF0000000000FFFF0000),
     .INIT_12(256'h000000E0F0381818000000070F1C1818181838F0E00000000C0C0C0C0C0C0C0C),
     .INIT_13(256'hC0C0C0C0C0C0FFFFC0E070381C0E070303070E1C3870E0C0FFFFC0C0C0C0C0C0),
     .INIT_14(256'h00081C3E7F7F7F3600FFFF0000000000003C7E7E7E7E3C00030303030303FFFF),
     .INIT_15(256'h003C7E66667E3C00C3E77E3C3C7EE7C318181C0F070000006060606060606060),
     .INIT_16(256'h181818FFFF18181800081C3E7F3E1C080606060606060606003C181866661818),
     .INIT_17(256'h0103070F1F3F7FFF003636763E03000018181818181818183030C0C03030C0C0),
     .INIT_18(256'h00000000000000FFFFFFFFFF00000000F0F0F0F0F0F0F0F00000000000000000),
     .INIT_19(256'h03030303030303033333CCCC3333CCCCC0C0C0C0C0C0C0C0FF00000000000000),
     .INIT_1A(256'h1818181F1F181818030303030303030380C0E0F0F8FCFEFF3333CCCC00000000),
     .INIT_1B(256'hFFFF000000000000181818F8F80000000000001F1F1818180F0F0F0F00000000),
     .INIT_1C(256'h181818F8F8181818181818FFFF000000000000FFFF1818181818181F1F000000),
     .INIT_1D(256'h000000000000FFFF0707070707070707E0E0E0E0E0E0E0E0C0C0C0C0C0C0C0C0),
     .INIT_1E(256'hF0F0F0F000000000FFFF030303030303FFFFFF00000000000000000000FFFFFF),
     .INIT_1F(256'h0F0F0F0FF0F0F0F000000000F0F0F0F0000000F8F8181818000000000F0F0F0F),
     .INIT_20(256'hFFC3999F9F9F99C3FF83999983999983FF9999998199C3E7FFC3999F919199C3),
     .INIT_21(256'hFFC39999919F99C3FF9F9F9F879F9F81FF819F9F879F9F81FF87939999999387),
     .INIT_22(256'hFF9993878F879399FFC793F3F3F3F3E1FFC3E7E7E7E7E7C3FF99999981999999),
     .INIT_23(256'hFFC39999999999C3FF99999181818999FF9C9C9C9480889CFF819F9F9F9F9F9F),
     .INIT_24(256'hFFC399F9C39F99C3FF99938783999983FFF1C399999999C3FF9F9F9F83999983),
     .INIT_25(256'hFF9C8880949C9C9CFFE7C39999999999FFC3999999999999FFE7E7E7E7E7E781),
     .INIT_26(256'hFFC3CFCFCFCFCFC3FF819FCFE7F3F981FFE7E7E7C3999999FF9999C3E7C39999),
     .INIT_27(256'hFFEFCF8080CFEFFFE7E7E7E781C3E7FFFFC3F3F3F3F3F3C3FF039DCF83CFEDF3),
     .INIT_28(256'hFF99990099009999FFFFFFFFFF999999FFE7FFFFE7E7E7E7FFFFFFFFFFFFFFFF),
     .INIT_29(256'hFFFFFFFFFFE7F3F9FFC09998C7C399C3FFB999CFE7F3999DFFE783F9C39FC1E7),
     .INIT_2A(256'hFFFFE7E781E7E7FFFFFF99C300C399FFFFCFE7F3F3F3E7CFFFF3E7CFCFCFE7F3),
     .INIT_2B(256'hFF9FCFE7F3F9FCFFFFE7E7FFFFFFFFFFFFFFFFFF81FFFFFFCFE7E7FFFFFFFFFF),
     .INIT_2C(256'hFFC399F9E3F999C3FF819FCFF3F999C3FF81E7E7E7C7E7E7FFC39999899199C3),
     .INIT_2D(256'hFFE7E7E7E7F39981FFC39999839F99C3FFC399F9F9839F81FFF9F98099E1F1F9),
     .INIT_2E(256'hCFE7E7FFFFE7FFFFFFFFE7FFFFE7FFFFFFC399F9C19999C3FFC39999C39999C3),
     .INIT_2F(256'hFFE7FFE7F3F999C3FF8FE7F3F9F3E78FFFFFFF81FF81FFFFFFF1E7CF9FCFE7F1),
     .INIT_30(256'hFFFFFF0000FFFFFFE7E7E7E7E7E7E7E7FFC1E38080C1E3F7FFFFFF0000FFFFFF),
     .INIT_31(256'hCFCFCFCFCFCFCFCFFFFF0000FFFFFFFFFFFFFFFFFF0000FFFFFFFFFF0000FFFF),
     .INIT_32(256'hFFFFFF1F0FC7E7E7FFFFFFF8F0E3E7E7E7E7C70F1FFFFFFFF3F3F3F3F3F3F3F3),
     .INIT_33(256'h3F3F3F3F3F3F00003F1F8FC7E3F1F8FCFCF8F1E3C78F1F3F00003F3F3F3F3F3F),
     .INIT_34(256'hFFF7E3C1808080C9FF0000FFFFFFFFFFFFC381818181C3FFFCFCFCFCFCFC0000),
     .INIT_35(256'hFFC381999981C3FF3C1881C3C381183CE7E7E3F0F8FFFFFF9F9F9F9F9F9F9F9F),
     .INIT_36(256'hE7E7E70000E7E7E7FFF7E3C180C1E3F7F9F9F9F9F9F9F9F9FFC3E7E79999E7E7),
     .INIT_37(256'hFEFCF8F0E0C08000FFC9C989C1FCFFFFE7E7E7E7E7E7E7E7CFCF3F3FCFCF3F3F),
     .INIT_38(256'hFFFFFFFFFFFFFF0000000000FFFFFFFF0F0F0F0F0F0F0F0FFFFFFFFFFFFFFFFF),
     .INIT_39(256'hFCFCFCFCFCFCFCFCCCCC3333CCCC33333F3F3F3F3F3F3F3F00FFFFFFFFFFFFFF),
     .INIT_3A(256'hE7E7E7E0E0E7E7E7FCFCFCFCFCFCFCFC7F3F1F0F07030100CCCC3333FFFFFFFF),
     .INIT_3B(256'h0000FFFFFFFFFFFFE7E7E70707FFFFFFFFFFFFE0E0E7E7E7F0F0F0F0FFFFFFFF),
     .INIT_3C(256'hE7E7E70707E7E7E7E7E7E70000FFFFFFFFFFFF0000E7E7E7E7E7E7E0E0FFFFFF),
     .INIT_3D(256'hFFFFFFFFFFFF0000F8F8F8F8F8F8F8F81F1F1F1F1F1F1F1F3F3F3F3F3F3F3F3F),
     .INIT_3E(256'h0F0F0F0FFFFFFFFF0000FCFCFCFCFCFC000000FFFFFFFFFFFFFFFFFFFF000000),
     .INIT_3F(256'hF0F0F0F00F0F0F0FFFFFFFFF0F0F0F0FFFFFFF0707E7E7E7FFFFFFFFF0F0F0F0),
     .INIT_40(256'h003C6060603C0000007C66667C606000003E663E063C0000003C62606E6E663C),
     .INIT_41(256'h7C063E66663E0000001818183E180E00003C607E663C0000003E66663E060600),
     .INIT_42(256'h00666C786C6060003C06060606000600003C181838001800006666667C606000),
     .INIT_43(256'h003C6666663C000000666666667C000000636B7F7F660000003C181818183800),
     .INIT_44(256'h007C063C603E000000606060667C000006063E66663E000060607C66667C0000),
     .INIT_45(256'h00363E7F6B63000000183C6666660000003E666666660000000E1818187E1800),
     .INIT_46(256'h003C30303030303C007E30180C7E0000780C3E666666000000663C183C660000),
     .INIT_47(256'h0010307F7F301000181818187E3C1800003C0C0C0C0C0C3C00FC62307C30120C),
     .INIT_48(256'h006666FF66FF6666000000000066666600180000181818180000000000000000),
     .INIT_49(256'h0000000000180C06003F6667383C663C00466630180C666200187C063C603E18),
     .INIT_4A(256'h000018187E1818000000663CFF3C66000030180C0C0C1830000C18303030180C),
     .INIT_4B(256'h006030180C0603000018180000000000000000007E0000003018180000000000),
     .INIT_4C(256'h003C66061C06663C007E60300C06663C007E181818381818003C6666766E663C),
     .INIT_4D(256'h00181818180C667E003C66667C60663C003C6606067C607E0006067F661E0E06),
     .INIT_4E(256'h30181800001800000000180000180000003C66063E66663C003C66663C66663C),
     .INIT_4F(256'h001800180C06663C0070180C060C18700000007E007E0000000E18306030180E),
     .INIT_50(256'h003C66606060663C007C66667C66667C006666667E663C18000000FFFF000000),
     .INIT_51(256'h003C66666E60663C006060607860607E007E60607860607E00786C6666666C78),
     .INIT_52(256'h00666C7870786C6600386C0C0C0C0C1E003C18181818183C006666667E666666),
     .INIT_53(256'h003C66666666663C0066666E7E7E7666006363636B7F7763007E606060606060),
     .INIT_54(256'h003C66063C60663C00666C787C66667C000E3C666666663C006060607C66667C),
     .INIT_55(256'h0063777F6B63636300183C6666666666003C666666666666001818181818187E),
     .INIT_56(256'h181818FFFF181818007E6030180C067E001818183C6666660066663C183C6666),
     .INIT_57(256'h66CC993366CC9933CCCC3333CCCC333318181818181818183030C0C03030C0C0),
     .INIT_58(256'h00000000000000FFFFFFFFFF00000000F0F0F0F0F0F0F0F00000000000000000),
     .INIT_59(256'h03030303030303033333CCCC3333CCCCC0C0C0C0C0C0C0C0FF00000000000000),
     .INIT_5A(256'h1818181F1F1818180303030303030303663399CC663399CC3333CCCC00000000),
     .INIT_5B(256'hFFFF000000000000181818F8F80000000000001F1F1818180F0F0F0F00000000),
     .INIT_5C(256'h181818F8F8181818181818FFFF000000000000FFFF1818181818181F1F000000),
     .INIT_5D(256'h000000000000FFFF0707070707070707E0E0E0E0E0E0E0E0C0C0C0C0C0C0C0C0),
     .INIT_5E(256'hF0F0F0F000000000006070786C060301FFFFFF00000000000000000000FFFFFF),
     .INIT_5F(256'h0F0F0F0FF0F0F0F000000000F0F0F0F0000000F8F8181818000000000F0F0F0F),
     .INIT_60(256'hFFC39F9F9FC3FFFFFF839999839F9FFFFFC199C1F9C3FFFFFFC3999F919199C3),
     .INIT_61(256'h83F9C19999C1FFFFFFE7E7E7C1E7F1FFFFC39F8199C3FFFFFFC19999C1F9F9FF),
     .INIT_62(256'hFF999387939F9FFFC3F9F9F9F9FFF9FFFFC3E7E7C7FFE7FFFF999999839F9FFF),
     .INIT_63(256'hFFC3999999C3FFFFFF9999999983FFFFFF9C94808099FFFFFFC3E7E7E7E7C7FF),
     .INIT_64(256'hFF83F9C39FC1FFFFFF9F9F9F9983FFFFF9F9C19999C1FFFF9F9F83999983FFFF),
     .INIT_65(256'hFFC9C180949CFFFFFFE7C3999999FFFFFFC199999999FFFFFFF1E7E7E781E7FF),
     .INIT_66(256'hFFC3CFCFCFCFCFC3FF81CFE7F381FFFF87F3C1999999FFFFFF99C3E7C399FFFF),
     .INIT_67(256'hFFEFCF8080CFEFFFE7E7E7E781C3E7FFFFC3F3F3F3F3F3C3FF039DCF83CFEDF3),
     .INIT_68(256'hFF99990099009999FFFFFFFFFF999999FFE7FFFFE7E7E7E7FFFFFFFFFFFFFFFF),
     .INIT_69(256'hFFFFFFFFFFE7F3F9FFC09998C7C399C3FFB999CFE7F3999DFFE783F9C39FC1E7),
     .INIT_6A(256'hFFFFE7E781E7E7FFFFFF99C300C399FFFFCFE7F3F3F3E7CFFFF3E7CFCFCFE7F3),
     .INIT_6B(256'hFF9FCFE7F3F9FCFFFFE7E7FFFFFFFFFFFFFFFFFF81FFFFFFCFE7E7FFFFFFFFFF),
     .INIT_6C(256'hFFC399F9E3F999C3FF819FCFF3F999C3FF81E7E7E7C7E7E7FFC39999899199C3),
     .INIT_6D(256'hFFE7E7E7E7F39981FFC39999839F99C3FFC399F9F9839F81FFF9F98099E1F1F9),
     .INIT_6E(256'hCFE7E7FFFFE7FFFFFFFFE7FFFFE7FFFFFFC399F9C19999C3FFC39999C39999C3),
     .INIT_6F(256'hFFE7FFE7F3F999C3FF8FE7F3F9F3E78FFFFFFF81FF81FFFFFFF1E7CF9FCFE7F1),
     .INIT_70(256'hFFC3999F9F9F99C3FF83999983999983FF9999998199C3E7FFFFFF0000FFFFFF),
     .INIT_71(256'hFFC39999919F99C3FF9F9F9F879F9F81FF819F9F879F9F81FF87939999999387),
     .INIT_72(256'hFF9993878F879399FFC793F3F3F3F3E1FFC3E7E7E7E7E7C3FF99999981999999),
     .INIT_73(256'hFFC39999999999C3FF99999181818999FF9C9C9C9480889CFF819F9F9F9F9F9F),
     .INIT_74(256'hFFC399F9C39F99C3FF99938783999983FFF1C399999999C3FF9F9F9F83999983),
     .INIT_75(256'hFF9C8880949C9C9CFFE7C39999999999FFC3999999999999FFE7E7E7E7E7E781),
     .INIT_76(256'hE7E7E70000E7E7E7FF819FCFE7F3F981FFE7E7E7C3999999FF9999C3E7C39999),
     .INIT_77(256'h993366CC993366CC3333CCCC3333CCCCE7E7E7E7E7E7E7E7CFCF3F3FCFCF3F3F),
     .INIT_78(256'hFFFFFFFFFFFFFF0000000000FFFFFFFF0F0F0F0F0F0F0F0FFFFFFFFFFFFFFFFF),
     .INIT_79(256'hFCFCFCFCFCFCFCFCCCCC3333CCCC33333F3F3F3F3F3F3F3F00FFFFFFFFFFFFFF),
     .INIT_7A(256'hE7E7E7E0E0E7E7E7FCFCFCFCFCFCFCFC99CC663399CC6633CCCC3333FFFFFFFF),
     .INIT_7B(256'h0000FFFFFFFFFFFFE7E7E70707FFFFFFFFFFFFE0E0E7E7E7F0F0F0F0FFFFFFFF),
     .INIT_7C(256'hE7E7E70707E7E7E7E7E7E70000FFFFFFFFFFFF0000E7E7E7E7E7E7E0E0FFFFFF),
     .INIT_7D(256'hFFFFFFFFFFFF0000F8F8F8F8F8F8F8F81F1F1F1F1F1F1F1F3F3F3F3F3F3F3F3F),
     .INIT_7E(256'h0F0F0F0FFFFFFFFFFF9F8F8793F9FCFE000000FFFFFFFFFFFFFFFFFFFF000000),
     .INIT_7F(256'hF0F0F0F00F0F0F0FFFFFFFFF0F0F0F0FFFFFFF0707E7E7E7FFFFFFFFF0F0F0F0),
     
     // The next set of INITP_xx are for the parity bits
     .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
     
     // The next set of INIT_xx are valid when configured as 36Kb
     .INITP_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_0F(256'h0000000000000000000000000000000000000000000000000000000000000000)
  ) BRAM_SINGLE_MACRO_inst_BLOCK_0 (
     .DO(DATA_OUT_BLOCK_0),       // Output data, width defined by READ_WIDTH parameter
     .ADDR(addr[11:0]),   // Input address, width defined by read/write port depth
     .CLK(clk),     // 1-bit input clock
     .DI(0),       // Input data port, width defined by WRITE_WIDTH parameter
     .EN(1),       // 1-bit input RAM enable
     .REGCE(0), // 1-bit input output register enable
     .RST(0),     // 1-bit input reset
     .WE(8'h00)        // Input write enable, width defined by write port depth
  );


//===============================================================================================


//===============================================================================================
  
     
 
  assign DO = DATA_OUT_BLOCK_0;
    
endmodule
