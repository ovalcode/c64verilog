`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05.07.2017 15:35:00
// Design Name: 
// Module Name: test
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module rom_kernal(
  input clk,
  input [12:0] addr,
  output [7:0] DO
  );
  
  
  
  wire [7:0] DATA_OUT_BLOCK_0;
  wire [7:0] DATA_OUT_BLOCK_1;
  wire nc_wire;
  reg [7:0] combined_data_out;
  reg bit_12_store;

    BRAM_SINGLE_MACRO #(
     .BRAM_SIZE("36Kb"), // Target BRAM, "18Kb" or "36Kb" 
     .DEVICE("7SERIES"), // Target Device: "7SERIES" 
     .DO_REG(0), // Optional output register (0 or 1)
     .INIT(36'h000000000), // Initial values on output port
     .INIT_FILE ("NONE"),
     .WRITE_WIDTH(8), // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
     .READ_WIDTH(8),  // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
     .SRVAL(36'h000000000), // Set/Reset value for port output
     .WRITE_MODE("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE" 
     .INIT_00(256'h69B505A24801E938F3F081691807A5BCCC20BAD420039088C961A5BC0F205685),
     .INIT_01(256'h20686F8500A9E05920BFA0C4A9BFB420B85320708556A5F510CA6994619561B4),
     .INIT_02(256'hBBC72072847185BA284C00A057A9E05D20BA282057A9BBCA207284718560BAB9),
     .INIT_03(256'h847185C8019005691872A471A5BA282072A4718572E602D098C871A4678571B1),
     .INIT_04(256'hF32020D03730BC2B200046B12868007A44359860E4D067C600A05CA9B8672072),
     .INIT_05(256'h8BA9E0E34C658522B1C8638522B108A0648522B1C8628522B104A023842286FF),
     .INIT_06(256'h8564A563A66286658562A565A6B86720E0A092A9BA2820E0A08DA9BBA22000A0),
     .INIT_07(256'h86388407D0F0C9BBD44C00A08BA2B8D720618580A9708561A5668500A9648663),
     .INIT_08(256'hC62060DCB0E4AD2060E2B0FFCF2060E8B0FFD220A4374C1EA202D0AAA6634C37),
     .INIT_09(256'h030DAE030CAD48030FAD4846A948E1A9B7F720AD8A2060D0B0FFE42060D6B0FF),
     .INIT_0A(256'h202BA92EA42DA6E1D42060030F8D68030E8C030D8E030C8D0800146C28030EAC),
     .INIT_0B(256'h1CA217F00AA557B0FFD5202CA42BA60AA5E1D4200A8500A92C01A96095B0FFD8),
     .INIT_0C(256'h374C1DA205F0BF29FFB72060AB1E4CA3A064A907F002C97AA517D01029FFB720),
     .INIT_0D(256'h1920A6774CA53320A68E20A52A4CAB1E20A3A076A92E842D860ED002C97BA5A4),
     .INIT_0E(256'hFFBA2000A001A2FFBD2000A9E0F94CC390FFC32049A5E21920600BB0FFC020E2),
     .INIT_0F(256'hFFBA4C49A6A88AE20020E20620FFBA20498600A0E20020E20620E25720E20620),
     .INIT_10(256'h1120FFBD2000A9AF084CF7D0007920AEFD2060686802D0007920B79E4CE20E20),
     .INIT_11(256'h2088019003E049A500A04A86E20020E20620FFBA2000A001A28A4986B79E20E2),
     .INIT_12(256'hA422A6B6A320AD9E20E20E20E20620FFBA2049A54AA6A88AE20020E20620FFBA),
     .INIT_13(256'h8500A9BCCC20BC0C20BB07206EA6E2A0E5A9BC0C20B86720E2A0E0A9FFBD4C23),
     .INIT_14(256'hBFB4201285FF4912A5093066A5B849200D104866A5B85020E2A0EAA9B853206F),
     .INIT_15(256'h4EA2E26B20128500A9BBCA20E0434CE2A0EFA9BFB420031068B86720E2A0EAA9),
     .INIT_16(256'hE29D4C48BB0F4C00A04EA9E2DC2012A5668500A9BBA22000A057A9E0F62000A0),
     .INIT_17(256'h870189689987F8FB0728861B2D1AE68405000000007FA2DA0F4983A2DA0F4981),
     .INIT_18(256'hA0BCA9079081C94861A5BFB42003104866A5A2DA0F498328E75DA586E1DF3523),
     .INIT_19(256'h760B60BFB44C031068B85020E2A0E0A9079081C968E04320E3A03EA9BB0F20B9),
     .INIT_1A(256'hEAB77D4C7064147DC1CB53DE7CCA671F0C7C10B0FC837BF5A6F41E79D3BD83B3),
     .INIT_1B(256'h00A9FFCC20000000008113AAAAAA7FC791CC4C7E3A9944927E7E8830637D7A51),
     .INIT_1C(256'h9AFBA2E42220E3BF20E45320A4744CA43A4C03308A03006C80A258A67A201385),
     .INIT_1D(256'hA95852C74F8060D0E93830E938EFF020C90AB03AC9EA60AD7BE602D07AE6E4D0),
     .INIT_1E(256'h04840385B1A0AAA906840585B3A091A903128C03118DB2A048A903108D54854C),
     .INIT_1F(256'h19A201FC8E01FD8E01A218851385688500A9538503A9F810CA7395E3A2BD1CA2),
     .INIT_20(256'hE602D02BE62B919800A03484338638843786FF9920382C842B86FF9C20381686),
     .INIT_21(256'hA060A9BDCD202CE538A5AA2BE53837A5AB1E20E4A073A9A408202CA42BA5602C),
     .INIT_22(256'h0060F710CA03009DE447BD0BA2AE86A7E4A71AA57CA483E38BA6444CAB1E20E4),
     .INIT_23(256'h4F43202A2A2A2A202020200D93000D4545524620534554594220434953414220),
     .INIT_24(256'h52204B3436200D0D2A2A2A2A2032562043495341422034362045524F444F4D4D),
     .INIT_25(256'hAAAAAAAAAAAAAAAAAA608A019068AAFFC92048810020204D4554535953204D41),
     .INIT_26(256'h60F3910286AD60AB8501A9A985AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA),
     .INIT_27(256'h006900AE013702D106060C700DE8111A1944261960F7D0A1C504D0C891A40269),
     .INIT_28(256'h02918D00A9E5A02060D3A4D6A6E56C20D384D68607B06019A028A260DCA000A2),
     .INIT_29(256'h0CA9028B8D04A902868D0EA9028C8D02898D0AA902908DEBA9028F8D48A9CF85),
     .INIT_2A(256'h18A2D995FFA9F3D01AE0E8C80190286918D994AA00A9A880090288ADCC85CD85),
     .INIT_2B(256'hA9E9F020F410CAD3852869180830D9B4D3A5D6A6D684D38400A0FA10CAE9FF20),
     .INIT_2C(256'hE5664CE5A020EA60E6ED4C03F0C9E4EA244CD585F610E82869180630D9B4E827),
     .INIT_2D(256'hE802779D0278BD00A20277AC60F7D0CACFFF9DECB8BD2FA2998500A99A8503A9),
     .INIT_2E(256'h0287AECEA50CF0CFA578F7F002928DCC85C6A5E7162060185898C6C6F5D0C6E4),
     .INIT_2F(256'h0DC9CFF0F7D0CA02769DECE6BDC6867809A210D083C9E5B420EA1320CF8400A0),
     .INIT_30(256'hA61B30C9A5D484D38402928C00A0C884C8F7D08803D020C9D1B1D084D5A4C8D0),
     .INIT_31(256'hD785D1B1D3A493F0D0A5488A48982BB00A90C8C5D385CAA512D0C9E4E59120D6),
     .INIT_32(256'h8500A917D0C8C4E68420D3E64009027004D0D4A6049080090210D724D7063F29),
     .INIT_33(256'h02D0DEC9D7A5A868AA68D7850DA9E7162003F003E09AA606F003E099A60DA9D0),
     .INIT_34(256'hAED8C602F0D8A6800902F0C7A640096022A9D4850149D4A508D022C96018FFA9),
     .INIT_35(256'hB0D3C5D5A5D3E6E8B32060581868AA68D44602F0D8A5A868E6B620EA13200286),
     .INIT_36(256'hB5E8D956D916D6A6D6C6E8EA20079019E0D6A6E9674C03F00292AD32F04FC93F),
     .INIT_37(256'hD38500A9E87C20D6C6E9F04CF9D0CA0330D9B5D585286918D5A5CAD9958009D9),
     .INIT_38(256'h8500A94898488AD7854860D384D5A4E56C20D686CA9DD06868D38606D0D6A660),
     .INIT_39(256'h203F2902D0DF29049060C9109020C9E8914C03D00DC9E7D44C0310D7A5D3A4D0),
     .INIT_3A(256'h20D38488E8A120E7734CE7012006D0982ED014C9E6974C03F0D8A6E6934CE684),
     .INIT_3B(256'hD4A64D10F3910286ADD19120A9EFD0D5C4C8F39188F3B1C8D19188D1B1C8EA24),
     .INIT_3C(256'h90D5C488D384E8B320C817D01DC9E5662003D013C9C78502D012C9E6974C03F0),
     .INIT_3D(256'hD6C6EAF0EC90D5C5D6E6A8286998181DD011C9E6A84CD38400A0E87C20D6C609),
     .INIT_3E(256'h039020C95EA902D07FC97F29EC444CE8CB20E6A84CE87C20F8D0D385049028E9),
     .INIT_3F(256'h4FC007D0D3C404D020C9D1B1D5A437D014C93FD0D4A6E8914C03D00DC9E6914C),
     .INIT_40(256'hADD19120A9EFD0D3C488F391C8F3B188D191C8D1B188EA2420D5A4E9652024F0),
     .INIT_41(256'hE938D3A5D6C637F0D6A616D011C9E6974C400905F0D8A6E6A84CD8E6F3910286),
     .INIT_42(256'h8488E8A12009F09812D01DC9C78500A904D012C925D0E56C202A10D385049028),
     .INIT_43(256'hD6A6C946EC4F4CE8CB208009E6A84CE5442006D013C9E6A84CE70120E6A84CD3),
     .INIT_44(256'hA84CE87C20D386D486C786D88600A2E56C4CD686F410D9B5E8EA2003D019E0E8),
     .INIT_45(256'hD0CA28691807F0D3C527A902A260D6C660F6D0CA28691807F0D3C500A902A2E6),
     .INIT_46(256'h1E9C9F1C05906002868E60F810CA04F0E8DADD0FA260D6E602F019E0D6A660F6),
     .INIT_47(256'hE802A5CEC9C6D6C6FFA248AFA548AEA548ADA548ACA59B9A9998979695819E1F),
     .INIT_48(256'h0210DAB47F29D9B500A2E9FF20EC30E9C820DAB5AC85ECF1BD0CB018E0E9F020),
     .INIT_49(256'hDC01ADDC008D7FA902A5EED6E6C310D9A5F1858009F1A5EFD018E0E8D9958009),
     .INIT_4A(256'h8568AE8568AF8568D6A6C684F9D088FCD0CAEA00A00BD028DC008D7FA908FBC9),
     .INIT_4B(256'hDA4CD6C6CA02A5AEE8EA200C900EF018E002A58EFB10D9B5E8D6A660AC8568AD),
     .INIT_4C(256'hB5AC85ECEFBD0CF00E9002A5ECE9F020CA19A248AFA548AEA548ADA548ACA5E6),
     .INIT_4D(256'hAEECD0CADA9580090210D9B47F29DAB50F9002A5EC17A2E9FF20E930E9C820D8),
     .INIT_4E(256'h60F51088F391AEB1D191ACB127A0E9E020AD8502880D0329E9584CE6DA2002A5),
     .INIT_4F(256'hA060D28502880D0329D9B5D185ECF0BD60AF85D8090329ADA5AE85ACA5EA2420),
     .INIT_50(256'hD191D3A498EA2420CD8502A9A8EA60F61088D19120A9E4DA20EA2420E9F02027),
     .INIT_51(256'hCD8514A925D0CDC629D0CCA5FFEA2060F485D8090329D2A5F385D1A560F3918A),
     .INIT_52(256'h1C208049CEA50286AE02878DF3B1EA2420CE85CFE611B0D1B10287AECF46D3A4),
     .INIT_53(256'h0DADEA872001851F2901A506D0C0A508D0200901A5C08400A00AF0102901A5EA),
     .INIT_54(256'hA9F58581A9A861F0FFE0DC01AEDC008DCB8440A0028D8D00A94068AA68A868DC),
     .INIT_55(256'hF003C90CB005C9F5B14816B04AF8D0DC01CDDC01AD4808A2DC008DFEA9F685EB),
     .INIT_56(256'h028F6C68CCD0DC008D2A6838DFD0CA0BB041C0C868CB840210028D8D028D0D08),
     .INIT_57(256'hF014C929F07FC949701630028A2C7F2936D0028C8C10A007F0C5C4AAF5B1CBA4),
     .INIT_58(256'h8B8C04A026D0028BCE2BD0028CCE05F0028CAC35D011C904F01DC908F020C90C),
     .INIT_59(256'hE802779D06B00289ECC6A68A0EF0FFE0028E8C028DACC584CBA41C1088C6A402),
     .INIT_5A(256'h188D0249D018AD1D300291ADEEF0028ECD15D003C9028DAD60DC008D7FA9C686),
     .INIT_5B(256'h78EC03EBC2EB81EAE04CF685EB7ABDF585EB79BDAA06A9029008C90AEB764CD0),
     .INIT_5C(256'h5548423847593758544643364452350145535A3441573311878685881D0D14EC),
     .INIT_5D(256'h51022032045F312F5E3D01133B2A5C2C403A2E2D4C502B4E4F4B4D304A493956),
     .INIT_5E(256'hC8C228C7D927D8D4C6C326C4D22501C5D3DA24C1D723918B8A898C9D8D94FF03),
     .INIT_5F(256'h02A022045F213FDE3D01935DC0A93CBA5B3EDDCCD0DBCECFCBCD30CAC929D6D5),
     .INIT_60(256'hBF9BA5B79ABDA3BBBC99ACB29801B1AEAD97B0B396918B8A898C9D8D94FF83D1),
     .INIT_61(256'hA095045F813FDE3D01935DDFA83CA45B3EDCB6AFA6AAB9A1A730B5A229BEB8B4),
     .INIT_62(256'h08C9E6A84CD0188DFD29D018AD0BD08EC909D00209D018AD07D00EC9FF83AB02),
     .INIT_63(256'hFFFFFFFFFFFFFFFFE6A84C02918D02912D7FA9EED009C9093002910D80A907D0),
     .INIT_64(256'h0E0F0B0D920A0912161508029E07191F181406031E04129CFF05131A9F01171C),
     .INIT_65(256'h00000000000000FFFF11FFFF05FF0690FF1E1FFFFF1DFF1CFF001BFFFF0C10FF),
     .INIT_66(256'h0004030201060E0000000000000F140008000000379B00000000000000000000),
     .INIT_67(256'h583008E0B890684018F0C8A0785028000D4E55520D44414F4C07060504030201),
     .INIT_68(256'hA3469446ED4020A366380A10942448F0A42020092C4009C098704820F8D0A880),
     .INIT_69(256'hEEB320EE9720EE8E2078DD008D0809DD00ADEE852003D03FC9EE972078958568),
     .INIT_6A(256'h20FB90EEA920FBB0EEA920FB90EEA9200A10A324EE852064B0EEA920EE972078),
     .INIT_6B(256'hEE8520EE972003D0EEA02005B095663F900AF8D0DD00CDDD00ADA58508A9EE8E),
     .INIT_6C(256'hADDC0DADDC0F8D19A9DC078D04A9D4D0A5C6DD008D1009DF29DD00ADEAEAEAEA),
     .INIT_6D(256'h00ADED362095854A901858FE1C2003A92C80A96058F4B0EEA9200AD00229DC0D),
     .INIT_6E(256'h3094246058FB30EEA920EE8520EDBE20EEA02078ED3620958560DD008DF729DD),
     .INIT_6F(256'h3FA92C5FA9DD008D0809DD00ADEE8E20786018958568ED40204805D094663805),
     .INIT_70(256'hFB10EEA920EE8520A58500A978EE974CEE8520AAFDD0CA0AA28AEDBE20ED1120),
     .INIT_71(256'hA5A51810F430EEA92007D00229DC0DADDC0DADEE9720DC0F8D19A9DC078D01A9),
     .INIT_72(256'hDD00CDDD00ADA58508A9CAD0A5E6FE1C2040A9EE8520EEA020EDB24C02A905F0),
     .INIT_73(256'hEE062003509024EEA020E4D0A5C6F5300AF8D0DD00CDDD00ADA466F5100AF8D0),
     .INIT_74(256'h60DD008DDF29DD00AD60DD008D1009DD00AD60DD008DEF29DD00AD601858A4A5),
     .INIT_75(256'h3047F0B4A560AAFDD0CAB8A28A600AF8D0DD00CDDD00AD60DD008D2009DD00AD),
     .INIT_76(256'h1C3014F002942C20A960B58504298A06F0B4C6BD85BD458ACA019000A2B6463F),
     .INIT_77(256'hE650E970EAD0EDF0BDA5F0D0B4E6DFD0B4C6E3100293ADB4C6CA01D0BDA51470),
     .INIT_78(256'h9DACB4860298AEB585BD8500A91E501D10DD012C07904A0294ADCBD0FFA2B4E6),
     .INIT_79(256'hA14DDD0D8D01A902978D02970D10A92C40A960029DEEB685F9B113F0029ECC02),
     .INIT_7A(256'hF0A8C633D0A9A660CACA0250CA01F002932C20A909A260DD0D8D02A18D800902),
     .INIT_7B(256'h90A9EFD0A86501A90A0293AD67F0A7A5A8C660AA66A746AB85AB45A7A50D3036),
     .INIT_7C(256'h2AF0029CCCC8029BACE4D34CEAD0A7A5EF3B4C02A9A98502A18D02A10DDD0D8D),
     .INIT_7D(256'hAB45A7A5B130B4F002942C20A9F791F8D0E84A04F009E00298AEAAA588029B8C),
     .INIT_7E(256'hF0F1D0AAA5EF7E4C02978D02970D02A92C80A92C04A92C01A9A6502CA97003F0),
     .INIT_7F(256'h01ADFB70DD012CF9D0022902A1AD20D01D10DD012C02A929904A0294AD9A85EC),
     
     // The next set of INITP_xx are for the parity bits
     .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
     
     // The next set of INIT_xx are valid when configured as 36Kb
     .INITP_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_0F(256'h0000000000000000000000000000000000000000000000000000000000000000)
  ) BRAM_SINGLE_MACRO_inst_BLOCK_0 (
     .DO(DATA_OUT_BLOCK_0),       // Output data, width defined by READ_WIDTH parameter
     .ADDR(addr[11:0]),   // Input address, width defined by read/write port depth
     .CLK(clk),     // 1-bit input clock
     .DI(0),       // Input data port, width defined by WRITE_WIDTH parameter
     .EN(1),       // 1-bit input RAM enable
     .REGCE(0), // 1-bit input output register enable
     .RST(0),     // 1-bit input reset
     .WE(8'h00)        // Input write enable, width defined by write port depth
  );


//===============================================================================================

  BRAM_SINGLE_MACRO #(
     .BRAM_SIZE("36Kb"), // Target BRAM, "18Kb" or "36Kb" 
     .DEVICE("7SERIES"), // Target Device: "7SERIES" 
     .DO_REG(0), // Optional output register (0 or 1)
     .INIT(36'h000000000), // Initial values on output port
     .INIT_FILE ("NONE"),
     .WRITE_WIDTH(8), // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
     .READ_WIDTH(8),  // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
     .SRVAL(36'h000000000), // Set/Reset value for port output
     .WRITE_MODE("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE" 
     .INIT_00(256'hF4F0029DCCC8029EACF02820601802978D40A9F9300770DD012CDD018D0209DD),
     .INIT_01(256'hA9DD058D029AADDD048D0299ADDD0E8D10A91EB04A02A1ADF9919EA588029E8C),
     .INIT_02(256'hAD10DD012C02A924F0082928904A0294AD998560DD0E8D11A9EF0620EF3B2081),
     .INIT_03(256'h02A1ADEF3B4C1890A9F9F00429DD01ADDD018DFD29DD01ADFAB04A02A1AD22F0),
     .INIT_04(256'h978D080960029CEEF7B102978DF7290BF0029BCC029CAC0297AD6018F3F01229),
     .INIT_05(256'h2F490D606802A18D00A9DD0D8D10A9F9D0032902A1AD11F002A1AD486000A902),
     .INIT_06(256'h502053534552500DA0524F46A0474E494843524145530DA320524F525245204F),
     .INIT_07(256'h4F2059414C5020262044524F434552205353455250C5504154204E4F2059414C),
     .INIT_08(256'hC74E495946495245560DA0474E495641530DC74E4944414F4C0DC5504154204E),
     .INIT_09(256'h99A56018F31028C8FFD2207F2908F0BDB90D109D248D4B4F0DA0444E554F460D),
     .INIT_0A(256'hA5CA85D3A50BD099A5601897A4F08620978418D002C9E5B44C780FF0C6A508D0),
     .INIT_0B(256'h16B0F1992097863FF002C938B0E6324CC885D5A5D08509D003C9E6324CC985D6),
     .INIT_0C(256'h41200BD0F80D206097A68A68AA606897A6A6C6FE1C2040A905D00DB0F1992048),
     .INIT_0D(256'hD000C9F7B0F14E20EE134C60180DA904F090A56018B2B1F0F0A68500A911B0F8),
     .INIT_0E(256'h8A9E85684AEDDD4C680490E7164C6804D003C99AA548EEF0E9D060290297ADF2),
     .INIT_0F(256'h68A86818B2919EA5A684C8B29100A002A90EB0F864200ED0F80D202390489848),
     .INIT_10(256'hF003C916F0BAA5F31F20F7014C03F0F30F20F1FC4CF017206000A902909EA5AA),
     .INIT_11(256'h200610B9A5ED0920AA60189985F70A4C03F060E0B9A6F04D4C03D002C914B012),
     .INIT_12(256'h4C03D0BAA5F31F20F7014C03F0F30F20F7074CE61090248AEDC720F2484CEDCC),
     .INIT_13(256'h10B9A5ED0C20AA60189A85EAF060E0B9A6EFE14C03D002C911B00FF003C9F70D),
     .INIT_14(256'hF0BAA5488AF31F20601802F0F31420F7074CE71090248AEDB92003D0EDBE2005),
     .INIT_15(256'hA9C801F0FAA5C801F0F8A5FE2720F48320F2F220681DD002C947B04CF003C950),
     .INIT_16(256'h6000A9680490F86420F1DD203800A9F7D02023F00F29B9A5F47D4CFA85F88500),
     .INIT_17(256'h599D0259B998A414F098E498C6AA68F64220F2F14CF76A2005A90BD062C9B9A5),
     .INIT_18(256'hBD60F8D00259DD1530CA98A68A908500A96018026D9D026DB902639D0263B902),
     .INIT_19(256'h03B099E4EDFE2003B09AE403A2988500A960B985026DBDBA850263BDB8850259),
     .INIT_1A(256'h4C03900AE098A6F6FE4C03D0F30F20F70A4C03D0B8A660998500A99A86EDEF20),
     .INIT_1B(256'h20059056F003C95AF002639DBAA5026D9DB9856009B9A502599DB8A598E6F6FB),
     .INIT_1C(256'hAF2036B0F817201FD00F29B9A5F7134C03B0F7D020F4094C03D002C94F90F3D5),
     .INIT_1D(256'h2004A917B0F83820F4B00C9020F0F72C20F7044C28F01890F7EA200AF0B7A5F5),
     .INIT_1E(256'h8500A9F6F0B7A4FA30B9A56018A68598B29102A900A007F060C0B9A4BFA9F76A),
     .INIT_1F(256'hDD20BBB100A00CF0B7A5F7074C6868051090A5EDB920F009B9A5ED0C20BAA590),
     .INIT_20(256'hEF4A20F2D004C0C8029399BBB10AF0B7C402978CF48320F6544CF6D0B7C4C8ED),
     .INIT_21(256'hE4EABDE4EBBCF4404CFEC0BDFEC1BC09D002A6ADAA0A1CF00F290293AD02988E),
     .INIT_22(256'h8D029BADF00D2003B00ADD01AD09904A0294ADFF2E200A0295AD02958D02968C),
     .INIT_23(256'hF0A938F986FA848805D0FAA5F786F8848805D0F8A5FE2720029D8D029EAD029C),
     .INIT_24(256'hC3866002A18C00A0DD008DDD000D04A9DD018DDD038D06A9DD0D8D7FA9FE2D4C),
     .INIT_25(256'hA6F7104C03D0B7A47B90F9F003C9F7134C03D0BAA5908500A9938503306CC484),
     .INIT_26(256'h50B04A4A90A5AE85EE1320EDC720B9A5ED0920BAA5F3D520B98560A9F5AF20B9),
     .INIT_27(256'h334C03D0FFE12090859025FDA9F5D220AF85C4A5AE85C3A508D08AAF85EE1320),
     .INIT_28(256'hAEE6AE912CFE1C2010A908F0AED100A00CF093A48AE8B04A4A90A5AAEE1320F6),
     .INIT_29(256'h134C03B0F7D020F7134C03B04AF7044C7990F64220EDEF20CB509024AFE602D0),
     .INIT_2A(256'h2990A5D3B053F0F72C20DAB05AF00B90F7EA2009F0B7A5F5AF2068B0F81720F7),
     .INIT_2B(256'hB103A0EFD0B9A504B0C485B2B1C8C385B2B101A0DDD003E011F001E04AD03810),
     .INIT_2C(256'hC4A5C185C3A5AF85C46598AE85C3658A18A8B2F102A0B2B104A0AAB2F101A0B2),
     .INIT_2D(256'h2F2017A015F0B7A5F12F200CA01E109DA560AFA4AEA61824F84A20F5D220C285),
     .INIT_2E(256'h84AE86F12B4C59A002F093A549A060F6D0B7C4C8FFD220BBB100A00CF0B7A4F1),
     .INIT_2F(256'hB7A4B98561A95F90F9F003C9F7134C03D0BAA503326CC28501B5C18500B5AAAF),
     .INIT_30(256'hA5EDDD20ACA5FB8E2000A0EDB920B9A5ED0C20BAA5F68F20F3D520F7104C03D0),
     .INIT_31(256'h20E5D0FCDB20603800A9F6422007D0FFE120EDDD20ACB116B0FCD120EDDD20AD),
     .INIT_32(256'h20F7134C03B04A6018EDFE20EDB920E009EF29B9A5ED0C20BAA51130B924EDFE),
     .INIT_33(256'hB0F8672012B0F76A208A01A202D00129B9A503A2F68F2025B0F838208D90F7D0),
     .INIT_34(256'hD0A2E600A2F5C14CF12F2051A0FB109DA5601824F76A2005A906F00229B9A50D),
     .INIT_35(256'hCDDC01ADA286A186A08606904FE9A0A51AE9A1A501E9A2A538A0E602D0A1E606),
     .INIT_36(256'hA2A57860918502D0E8DC008DF8D0DC01ECDC01AEDC008EBDA21330AAF8D0DC01),
     .INIT_37(256'h02A92C01A96028C685FFCC200807D07FC991A56058A084A186A28578A0A4A1A6),
     .INIT_38(256'h200A509D2400A0FFCC204809A92C08A92C07A92C06A92C05A92C04A92C03A92C),
     .INIT_39(256'hC92AF005C9B2B100A032B0938568F841204893A5603868FFD22030094868F12F),
     .INIT_3A(256'hD015C0C8FFD220B2B105A0F12F2063A017109D24AAE1D004C904F003C908F001),
     .INIT_3B(256'hA9BFA048AEA548AFA548C1A548C2A55E90F7D0209E85608818EAE4E020A1A5F6),
     .INIT_3C(256'h84C8B291AFA5C8B291AEA5C8B291C2A5C8B291C1A5C8B2919EA5FBD088B29120),
     .INIT_3D(256'h6B20AB8569A9F7D720EED09FE69EE6B2919FA4BBB10CF0B7C49EA49E8400A09F),
     .INIT_3E(256'hC06918C1858AF7D0206002C0B3A4B2A66098C28568C18568AF8568AE8568A8F8),
     .INIT_3F(256'hD19FA4BBB110F0B7C49E8400A09F8405A01DB0F72C2060AF850069C28598AE85),
     .INIT_40(256'h2F201BA01AF0F82E2060C0C0A6A4A6E6F7D0206018ECD09EA49FE69EE6E7D0B2),
     .INIT_41(256'hD02EA0F9F0F82E206018012402D0012410A9F12F4C6AA0F8D0F82E20F8D020F1),
     .INIT_42(256'h90A99C859F859E85B085B485AA8500A9781FB0F81720F7D7209385908500A9DD),
     .INIT_43(256'hDC0EADDC0D8DDC0D8C7FA008A282A9786CB0F83820AB8514A9F7D72011D00EA2),
     .INIT_44(256'hA08D0315AD029F8D0314ADD0118DEF29D011ADF0A42002A28D9129DC0F8D1909),
     .INIT_45(256'hA0AD58F8D0CAFDD088FFA0FFA2C08501851F2901A5FB9720BE8502A9FCBD2002),
     .INIT_46(256'hA08D00A9686838FC93200BD018FFE120F8BE4CF6BC20F8D02015F0180315CD02),
     .INIT_47(256'h06ADAA2AB1062AB1062A0130B02400A9B185B16518B065180A0AB0A5B1866002),
     .INIT_48(256'hF01029DC0DAD02A48DDC0E8D02A2ADDC058DDC076D8ADC048DB165F99016C9DC),
     .INIT_49(256'hDC068CAAB186F2D0DC07ECDC06ED98FFA0DC07AE6058FF434C482AA948F9A909),
     .INIT_4A(256'hB1C53C6918B0A5B1664AB1664AB186B1E59802A38DDC0DADDC0F8D19A9DC078C),
     .INIT_4B(256'h17B0B1C5B0652669E81CB0B1C5B065306900A21B30A3A6FA604C03F09CA64AB0),
     .INIT_4C(256'h9265B1E513E938A9C602B0A9E619D0A8851DF0B4A5FA104C0390B1C5B0652C69),
     .INIT_4D(256'hA48500A916D002A4AD05D0012902A3AD22F0B4A5D7862BF0A4850149A4A59285),
     .INIT_4E(256'hB0E62CB0C6033007F092A5FEBC4CB9D09BA5F8E220A6A2BF303010A3A502A48D),
     .INIT_4F(256'hD2F0B4A59B859B458AB5B09685B99010C9BD30A9A5A0D08A0FD0D7E4928500A9),
     .INIT_50(256'h46F9974C0330A3A507F0B4A504F096A5FEBC4CF8E220DAA2BF66D746C530A3C6),
     .INIT_51(256'h8D81A9968500A9A88526F096A511D0B4A59CE6F8E220AA0AB065B1E53893A9B1),
     .INIT_52(256'hFEBC4CB685A905A8A5BD85BFA5DC0D8D01A9B48500A909F0B58596A5B485DC0D),
     .INIT_53(256'hA90BD0CABEA60CD0B5A51710AA240FA9A78502F0BEA5F8E220DAA29C85FB9720),
     .INIT_54(256'h0330BDA54AA7A5F1D0B6A5F5D0B5A518D03170FEBC4CAA8500A904D0FE1C2008),
     .INIT_55(256'hCAD0AA8580A9D0F0AB8500A9FB8E20AA8540A9DDD0AAC6AA850F2915B0181890),
     .INIT_56(256'hA00CF093A52DF0CAA7A6FB484C0390FCD120FB4A4C00A9FE1C2004A90AF0B5A5),
     .INIT_57(256'h009DACA501019DADA59EA63E909EE43DA24BF0B6A5B68501A904F0ACD1BDA500),
     .INIT_58(256'h9FE69FE627D00101DDADA52ED00100DDACA535F09EE49FA6FB3A4C9E86E8E801),
     .INIT_59(256'hA5A805D093A509D0FE1C2010A907F0B6A5B684C817F0ACD100A0BDA50BF093A5),
     .INIT_5A(256'h08F0A7C6BE860230CABEA6DC0DAEDC0D8E01A278AA8580A943D0FCDB20AC91BD),
     .INIT_5B(256'hF290FCD120FCDB20AB85AB45ACB1AB8400A0FB8E20FC932023F0BE8527D09EA5),
     .INIT_5C(256'h85A48500A9A38508A960AC85C1A5AD85C2A5FEBC4CFE1C2020A905F0BD45ABA5),
     .INIT_5D(256'hA5DC0F8D19A9DC0DADDC078EDC068D00A2B0A9029060A94ABDA560A9859B85A8),
     .INIT_5E(256'h2910B6A5A8E62FD0FBB12001A210A912D0A8A53C30B666386008290185084901),
     .INIT_5F(256'h49BDA50FF0A4850149A4A514D0FBA62019D0A9E61DD0FBAD2009D0A9A5FC574C),
     .INIT_60(256'h00A212F0A5A558FB9720F3103AF0A3A5A3C6BD46FEBC4C9B859B450129BD8501),
     .INIT_61(256'hA0CAB0BD85D7A5ADE691D00A90FCD120D9D0BD85800902D002E0BEA6A5C6D786),
     .INIT_62(256'h50A9FCCA2003D0BEC6FEBC4CBD8501499BA5BBD0FCDB20D785D745BD85ACB100),
     .INIT_63(256'hBD200AA2D810ABC6FB9720DFD0A7C6E3D0FBAF2078A9EAD0FCBD207808A2A785),
     .INIT_64(256'hFCCA20D0118D1009D011AD780883D0B686A58609A2FB8E2030F0BEA5ABE658FC),
     .INIT_65(256'hFD93BD97F0FC9320602803148D029FAD03158D09F002A0ADFDDD20DC0D8D7FA9),
     .INIT_66(256'hE602D0ACE660AFE5ADA5AEE5ACA538600185200901A56003158DFD94BD03148D),
     .INIT_67(256'h6C58FF5B20FD1520FD5020FDA320D0168E80006C03D0FD0220D89A78FFA260AD),
     .INIT_68(256'h1FA0C484C38618FDA030A23038CDC2C360F5D0CA03D08003DDFD0FBD05A2A000),
     .INIT_69(256'hF333F250F20EF291F34AFE47FE66EA3160F11088031499C391C3B102B00314B9),
     .INIT_6A(256'hA2F4D0C8030099020099000299A800A9F5EDF4A5FE66F32FF13EF6EDF1CAF157),
     .INIT_6B(256'h08D0C1D1C1912A0FD0C1D1C19155A9AAC1B1C2E6C28503A9A8B384B28603A03C),
     .INIT_6C(256'h31FBCDFC6A6002888D04A902828D08A9FE2D2018C2A4AA98E4F0E8D0C8C1918A),
     .INIT_6D(256'h038E00A2DD0F8DDC0F8DDD0E8DDC0E8D08A9DC008DDD0D8DDC0D8D7FA9F92CEA),
     .INIT_6E(256'h02A6AD00852FA90185E7A9DD028D3FA9DD008D07A9DC028ECAD4188EDD038EDC),
     .INIT_6F(256'h60BC84BB86B785FF6E4CDC058D42A9DC048D95A9FDF34C40A9DC048D25A90AF0),
     .INIT_70(256'h9085900590A59D85606802978D00A9480297AD0DD002C9BAA560B984BA86B885),
     .INIT_71(256'h8C02818E0282AC0281AE06906002848C02838E0284AC0283AE06906002858D60),
     .INIT_72(256'hBC2080026C03D0FD02201C30DD0DACDD0D8D7FA94898488A4803186C78600282),
     .INIT_73(256'hFB29DD00AD28F00129AA02A12D98A0026CE51820FDA320FD15200CD0FFE120F6),
     .INIT_74(256'hEEBB20FF0720FE9D4CFED62006F002290DF012298ADD0D8D02A1ADDD008DB505),
     .INIT_75(256'hAA68A868DD0D8D02A1ADFF072003F010298AFEB64CFED62006F002298AFEB64C),
     .INIT_76(256'hDD06ADA7850129DD01AD007100B8014602F006450CED0E7411C51A3E27C14068),
     .INIT_77(256'h068DFFA9DD0D8D02A1ADDD0F8D11A9DD078D029A6DDD07ADDD068D02996D1CE9),
     .INIT_78(256'h02A18D02A14D12A9DD0F8D11A9DD078D0296ADDD068D0295ADEF594CDD078DDD),
     .INIT_79(256'h029A8D00699802998DC8698AA82A0296ADAA60A8860298AEDD078DDD068DFFA9),
     .INIT_7A(256'h12ADE5182003146C03166C03F010290104BDBA4898488A4848EF296808EAEA60),
     .INIT_7B(256'hEE8E4CDC0E8D11098029DC0EADDC0D8D81A9FDDD4C02A68D0129D019ADFBD0D0),
     .INIT_7C(256'h4CFE344CFE254CEDC74CEDB94CFE184CFD1A4CFD154CFD504CFDA34CFF5B4C03),
     .INIT_7D(256'hFDF94CFE004CFE074CED094CED0C4CEDFE4CEDEF4CEDDD4CEE134CFE214CEA87),
     .INIT_7E(256'hDD4CF6E44CF5DD4CF49E4C03266C03246C03226C03206C031E6C031C6C031A6C),
     .INIT_7F(256'hFF48FCE2FE4359425252E5004CE50A4CE5054CF69B4C032C6C032A6C03286CF6),
     
     // The next set of INITP_xx are for the parity bits
     .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
     
     // The next set of INIT_xx are valid when configured as 36Kb
     .INITP_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
     .INITP_0F(256'h0000000000000000000000000000000000000000000000000000000000000000)
  ) BRAM_SINGLE_MACRO_inst_BLOCK_3 (
     .DO(DATA_OUT_BLOCK_1),       // Output data, width defined by READ_WIDTH parameter
     .ADDR(addr[11:0]),   // Input address, width defined by read/write port depth
     .CLK(clk),     // 1-bit input clock
     .DI(0),       // Input data port, width defined by WRITE_WIDTH parameter
     .EN(1),       // 1-bit input RAM enable
     .REGCE(0), // 1-bit input output register enable
     .RST(0),     // 1-bit input reset
     .WE(8'h00)        // Input write enable, width defined by write port depth
  );


//===============================================================================================
  
  always @(posedge clk)
  bit_12_store <= addr[12];
     
  always @*
  case (bit_12_store)
    1'b0: combined_data_out = DATA_OUT_BLOCK_0;
    1'b1: combined_data_out = DATA_OUT_BLOCK_1;
    default:  combined_data_out = 0;
  endcase
 
  assign DO = combined_data_out;
  
    
endmodule
